`include "../packages.sv"

module reduce_angle
    import fixed_pkg::fixed_t;
(
    input fixed_t angle,
    output fixed_t reduced_angle
);

endmodule: reduce_angle
