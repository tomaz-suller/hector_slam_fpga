`include "../packages.sv"

module tangent_lut
    import fixed_pkg::fixed_t;
(
    input fixed_t in,
    output fixed_t out
);

endmodule: tangent_lut
