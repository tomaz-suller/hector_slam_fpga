module tangent_lut
(
    input logic [31:0] in,
    output logic [31:0] out
);

endmodule: tangent_lut
