module tangent_lut
(
    input logic [31:0] in,
    output logic [31:0] out
);

    logic [11:0] truncated_in;
    assign truncated_in = in [18:7];

    always_comb begin
        case (truncated_in)
            12'b000000000000: out = 32'b00000000000000000000000000000000;
            12'b000000000001: out = 32'b00000000000000000000000010000000;
            12'b000000000010: out = 32'b00000000000000000000000100000000;
            12'b000000000011: out = 32'b00000000000000000000000110000000;
            12'b000000000100: out = 32'b00000000000000000000001000000000;
            12'b000000000101: out = 32'b00000000000000000000001010000000;
            12'b000000000110: out = 32'b00000000000000000000001100000000;
            12'b000000000111: out = 32'b00000000000000000000001110000000;
            12'b000000001000: out = 32'b00000000000000000000010000000000;
            12'b000000001001: out = 32'b00000000000000000000010010000000;
            12'b000000001010: out = 32'b00000000000000000000010100000000;
            12'b000000001011: out = 32'b00000000000000000000010110000000;
            12'b000000001100: out = 32'b00000000000000000000011000000000;
            12'b000000001101: out = 32'b00000000000000000000011010000000;
            12'b000000001110: out = 32'b00000000000000000000011100000000;
            12'b000000001111: out = 32'b00000000000000000000011110000000;
            12'b000000010000: out = 32'b00000000000000000000100000000000;
            12'b000000010001: out = 32'b00000000000000000000100010000000;
            12'b000000010010: out = 32'b00000000000000000000100100000000;
            12'b000000010011: out = 32'b00000000000000000000100110000000;
            12'b000000010100: out = 32'b00000000000000000000101000000000;
            12'b000000010101: out = 32'b00000000000000000000101010000000;
            12'b000000010110: out = 32'b00000000000000000000101100000000;
            12'b000000010111: out = 32'b00000000000000000000101110000000;
            12'b000000011000: out = 32'b00000000000000000000110000000000;
            12'b000000011001: out = 32'b00000000000000000000110010000000;
            12'b000000011010: out = 32'b00000000000000000000110100000000;
            12'b000000011011: out = 32'b00000000000000000000110110000000;
            12'b000000011100: out = 32'b00000000000000000000111000000000;
            12'b000000011101: out = 32'b00000000000000000000111010000000;
            12'b000000011110: out = 32'b00000000000000000000111100000000;
            12'b000000011111: out = 32'b00000000000000000000111110000000;
            12'b000000100000: out = 32'b00000000000000000001000000000000;
            12'b000000100001: out = 32'b00000000000000000001000010000000;
            12'b000000100010: out = 32'b00000000000000000001000100000000;
            12'b000000100011: out = 32'b00000000000000000001000110000000;
            12'b000000100100: out = 32'b00000000000000000001001000000000;
            12'b000000100101: out = 32'b00000000000000000001001010000000;
            12'b000000100110: out = 32'b00000000000000000001001100000000;
            12'b000000100111: out = 32'b00000000000000000001001110000000;
            12'b000000101000: out = 32'b00000000000000000001010000000000;
            12'b000000101001: out = 32'b00000000000000000001010010000000;
            12'b000000101010: out = 32'b00000000000000000001010100000000;
            12'b000000101011: out = 32'b00000000000000000001010110000000;
            12'b000000101100: out = 32'b00000000000000000001011000000000;
            12'b000000101101: out = 32'b00000000000000000001011010000000;
            12'b000000101110: out = 32'b00000000000000000001011100000000;
            12'b000000101111: out = 32'b00000000000000000001011110000001;
            12'b000000110000: out = 32'b00000000000000000001100000000001;
            12'b000000110001: out = 32'b00000000000000000001100010000001;
            12'b000000110010: out = 32'b00000000000000000001100100000001;
            12'b000000110011: out = 32'b00000000000000000001100110000001;
            12'b000000110100: out = 32'b00000000000000000001101000000001;
            12'b000000110101: out = 32'b00000000000000000001101010000001;
            12'b000000110110: out = 32'b00000000000000000001101100000001;
            12'b000000110111: out = 32'b00000000000000000001101110000001;
            12'b000000111000: out = 32'b00000000000000000001110000000001;
            12'b000000111001: out = 32'b00000000000000000001110010000001;
            12'b000000111010: out = 32'b00000000000000000001110100000001;
            12'b000000111011: out = 32'b00000000000000000001110110000010;
            12'b000000111100: out = 32'b00000000000000000001111000000010;
            12'b000000111101: out = 32'b00000000000000000001111010000010;
            12'b000000111110: out = 32'b00000000000000000001111100000010;
            12'b000000111111: out = 32'b00000000000000000001111110000010;
            12'b000001000000: out = 32'b00000000000000000010000000000010;
            12'b000001000001: out = 32'b00000000000000000010000010000010;
            12'b000001000010: out = 32'b00000000000000000010000100000010;
            12'b000001000011: out = 32'b00000000000000000010000110000011;
            12'b000001000100: out = 32'b00000000000000000010001000000011;
            12'b000001000101: out = 32'b00000000000000000010001010000011;
            12'b000001000110: out = 32'b00000000000000000010001100000011;
            12'b000001000111: out = 32'b00000000000000000010001110000011;
            12'b000001001000: out = 32'b00000000000000000010010000000011;
            12'b000001001001: out = 32'b00000000000000000010010010000011;
            12'b000001001010: out = 32'b00000000000000000010010100000100;
            12'b000001001011: out = 32'b00000000000000000010010110000100;
            12'b000001001100: out = 32'b00000000000000000010011000000100;
            12'b000001001101: out = 32'b00000000000000000010011010000100;
            12'b000001001110: out = 32'b00000000000000000010011100000100;
            12'b000001001111: out = 32'b00000000000000000010011110000101;
            12'b000001010000: out = 32'b00000000000000000010100000000101;
            12'b000001010001: out = 32'b00000000000000000010100010000101;
            12'b000001010010: out = 32'b00000000000000000010100100000101;
            12'b000001010011: out = 32'b00000000000000000010100110000101;
            12'b000001010100: out = 32'b00000000000000000010101000000110;
            12'b000001010101: out = 32'b00000000000000000010101010000110;
            12'b000001010110: out = 32'b00000000000000000010101100000110;
            12'b000001010111: out = 32'b00000000000000000010101110000110;
            12'b000001011000: out = 32'b00000000000000000010110000000110;
            12'b000001011001: out = 32'b00000000000000000010110010000111;
            12'b000001011010: out = 32'b00000000000000000010110100000111;
            12'b000001011011: out = 32'b00000000000000000010110110000111;
            12'b000001011100: out = 32'b00000000000000000010111000000111;
            12'b000001011101: out = 32'b00000000000000000010111010001000;
            12'b000001011110: out = 32'b00000000000000000010111100001000;
            12'b000001011111: out = 32'b00000000000000000010111110001000;
            12'b000001100000: out = 32'b00000000000000000011000000001001;
            12'b000001100001: out = 32'b00000000000000000011000010001001;
            12'b000001100010: out = 32'b00000000000000000011000100001001;
            12'b000001100011: out = 32'b00000000000000000011000110001001;
            12'b000001100100: out = 32'b00000000000000000011001000001010;
            12'b000001100101: out = 32'b00000000000000000011001010001010;
            12'b000001100110: out = 32'b00000000000000000011001100001010;
            12'b000001100111: out = 32'b00000000000000000011001110001011;
            12'b000001101000: out = 32'b00000000000000000011010000001011;
            12'b000001101001: out = 32'b00000000000000000011010010001011;
            12'b000001101010: out = 32'b00000000000000000011010100001100;
            12'b000001101011: out = 32'b00000000000000000011010110001100;
            12'b000001101100: out = 32'b00000000000000000011011000001100;
            12'b000001101101: out = 32'b00000000000000000011011010001101;
            12'b000001101110: out = 32'b00000000000000000011011100001101;
            12'b000001101111: out = 32'b00000000000000000011011110001101;
            12'b000001110000: out = 32'b00000000000000000011100000001110;
            12'b000001110001: out = 32'b00000000000000000011100010001110;
            12'b000001110010: out = 32'b00000000000000000011100100001111;
            12'b000001110011: out = 32'b00000000000000000011100110001111;
            12'b000001110100: out = 32'b00000000000000000011101000001111;
            12'b000001110101: out = 32'b00000000000000000011101010010000;
            12'b000001110110: out = 32'b00000000000000000011101100010000;
            12'b000001110111: out = 32'b00000000000000000011101110010001;
            12'b000001111000: out = 32'b00000000000000000011110000010001;
            12'b000001111001: out = 32'b00000000000000000011110010010010;
            12'b000001111010: out = 32'b00000000000000000011110100010010;
            12'b000001111011: out = 32'b00000000000000000011110110010010;
            12'b000001111100: out = 32'b00000000000000000011111000010011;
            12'b000001111101: out = 32'b00000000000000000011111010010011;
            12'b000001111110: out = 32'b00000000000000000011111100010100;
            12'b000001111111: out = 32'b00000000000000000011111110010100;
            12'b000010000000: out = 32'b00000000000000000100000000010101;
            12'b000010000001: out = 32'b00000000000000000100000010010101;
            12'b000010000010: out = 32'b00000000000000000100000100010110;
            12'b000010000011: out = 32'b00000000000000000100000110010110;
            12'b000010000100: out = 32'b00000000000000000100001000010111;
            12'b000010000101: out = 32'b00000000000000000100001010010111;
            12'b000010000110: out = 32'b00000000000000000100001100011000;
            12'b000010000111: out = 32'b00000000000000000100001110011001;
            12'b000010001000: out = 32'b00000000000000000100010000011001;
            12'b000010001001: out = 32'b00000000000000000100010010011010;
            12'b000010001010: out = 32'b00000000000000000100010100011010;
            12'b000010001011: out = 32'b00000000000000000100010110011011;
            12'b000010001100: out = 32'b00000000000000000100011000011011;
            12'b000010001101: out = 32'b00000000000000000100011010011100;
            12'b000010001110: out = 32'b00000000000000000100011100011101;
            12'b000010001111: out = 32'b00000000000000000100011110011101;
            12'b000010010000: out = 32'b00000000000000000100100000011110;
            12'b000010010001: out = 32'b00000000000000000100100010011111;
            12'b000010010010: out = 32'b00000000000000000100100100011111;
            12'b000010010011: out = 32'b00000000000000000100100110100000;
            12'b000010010100: out = 32'b00000000000000000100101000100001;
            12'b000010010101: out = 32'b00000000000000000100101010100001;
            12'b000010010110: out = 32'b00000000000000000100101100100010;
            12'b000010010111: out = 32'b00000000000000000100101110100011;
            12'b000010011000: out = 32'b00000000000000000100110000100011;
            12'b000010011001: out = 32'b00000000000000000100110010100100;
            12'b000010011010: out = 32'b00000000000000000100110100100101;
            12'b000010011011: out = 32'b00000000000000000100110110100101;
            12'b000010011100: out = 32'b00000000000000000100111000100110;
            12'b000010011101: out = 32'b00000000000000000100111010100111;
            12'b000010011110: out = 32'b00000000000000000100111100101000;
            12'b000010011111: out = 32'b00000000000000000100111110101000;
            12'b000010100000: out = 32'b00000000000000000101000000101001;
            12'b000010100001: out = 32'b00000000000000000101000010101010;
            12'b000010100010: out = 32'b00000000000000000101000100101011;
            12'b000010100011: out = 32'b00000000000000000101000110101100;
            12'b000010100100: out = 32'b00000000000000000101001000101100;
            12'b000010100101: out = 32'b00000000000000000101001010101101;
            12'b000010100110: out = 32'b00000000000000000101001100101110;
            12'b000010100111: out = 32'b00000000000000000101001110101111;
            12'b000010101000: out = 32'b00000000000000000101010000110000;
            12'b000010101001: out = 32'b00000000000000000101010010110001;
            12'b000010101010: out = 32'b00000000000000000101010100110010;
            12'b000010101011: out = 32'b00000000000000000101010110110011;
            12'b000010101100: out = 32'b00000000000000000101011000110011;
            12'b000010101101: out = 32'b00000000000000000101011010110100;
            12'b000010101110: out = 32'b00000000000000000101011100110101;
            12'b000010101111: out = 32'b00000000000000000101011110110110;
            12'b000010110000: out = 32'b00000000000000000101100000110111;
            12'b000010110001: out = 32'b00000000000000000101100010111000;
            12'b000010110010: out = 32'b00000000000000000101100100111001;
            12'b000010110011: out = 32'b00000000000000000101100110111010;
            12'b000010110100: out = 32'b00000000000000000101101000111011;
            12'b000010110101: out = 32'b00000000000000000101101010111100;
            12'b000010110110: out = 32'b00000000000000000101101100111101;
            12'b000010110111: out = 32'b00000000000000000101101110111110;
            12'b000010111000: out = 32'b00000000000000000101110000111111;
            12'b000010111001: out = 32'b00000000000000000101110011000000;
            12'b000010111010: out = 32'b00000000000000000101110101000001;
            12'b000010111011: out = 32'b00000000000000000101110111000010;
            12'b000010111100: out = 32'b00000000000000000101111001000011;
            12'b000010111101: out = 32'b00000000000000000101111011000100;
            12'b000010111110: out = 32'b00000000000000000101111101000110;
            12'b000010111111: out = 32'b00000000000000000101111111000111;
            12'b000011000000: out = 32'b00000000000000000110000001001000;
            12'b000011000001: out = 32'b00000000000000000110000011001001;
            12'b000011000010: out = 32'b00000000000000000110000101001010;
            12'b000011000011: out = 32'b00000000000000000110000111001011;
            12'b000011000100: out = 32'b00000000000000000110001001001100;
            12'b000011000101: out = 32'b00000000000000000110001011001110;
            12'b000011000110: out = 32'b00000000000000000110001101001111;
            12'b000011000111: out = 32'b00000000000000000110001111010000;
            12'b000011001000: out = 32'b00000000000000000110010001010001;
            12'b000011001001: out = 32'b00000000000000000110010011010010;
            12'b000011001010: out = 32'b00000000000000000110010101010100;
            12'b000011001011: out = 32'b00000000000000000110010111010101;
            12'b000011001100: out = 32'b00000000000000000110011001010110;
            12'b000011001101: out = 32'b00000000000000000110011011010111;
            12'b000011001110: out = 32'b00000000000000000110011101011001;
            12'b000011001111: out = 32'b00000000000000000110011111011010;
            12'b000011010000: out = 32'b00000000000000000110100001011011;
            12'b000011010001: out = 32'b00000000000000000110100011011101;
            12'b000011010010: out = 32'b00000000000000000110100101011110;
            12'b000011010011: out = 32'b00000000000000000110100111011111;
            12'b000011010100: out = 32'b00000000000000000110101001100001;
            12'b000011010101: out = 32'b00000000000000000110101011100010;
            12'b000011010110: out = 32'b00000000000000000110101101100100;
            12'b000011010111: out = 32'b00000000000000000110101111100101;
            12'b000011011000: out = 32'b00000000000000000110110001100110;
            12'b000011011001: out = 32'b00000000000000000110110011101000;
            12'b000011011010: out = 32'b00000000000000000110110101101001;
            12'b000011011011: out = 32'b00000000000000000110110111101011;
            12'b000011011100: out = 32'b00000000000000000110111001101100;
            12'b000011011101: out = 32'b00000000000000000110111011101110;
            12'b000011011110: out = 32'b00000000000000000110111101101111;
            12'b000011011111: out = 32'b00000000000000000110111111110001;
            12'b000011100000: out = 32'b00000000000000000111000001110010;
            12'b000011100001: out = 32'b00000000000000000111000011110100;
            12'b000011100010: out = 32'b00000000000000000111000101110101;
            12'b000011100011: out = 32'b00000000000000000111000111110111;
            12'b000011100100: out = 32'b00000000000000000111001001111001;
            12'b000011100101: out = 32'b00000000000000000111001011111010;
            12'b000011100110: out = 32'b00000000000000000111001101111100;
            12'b000011100111: out = 32'b00000000000000000111001111111110;
            12'b000011101000: out = 32'b00000000000000000111010001111111;
            12'b000011101001: out = 32'b00000000000000000111010100000001;
            12'b000011101010: out = 32'b00000000000000000111010110000011;
            12'b000011101011: out = 32'b00000000000000000111011000000100;
            12'b000011101100: out = 32'b00000000000000000111011010000110;
            12'b000011101101: out = 32'b00000000000000000111011100001000;
            12'b000011101110: out = 32'b00000000000000000111011110001001;
            12'b000011101111: out = 32'b00000000000000000111100000001011;
            12'b000011110000: out = 32'b00000000000000000111100010001101;
            12'b000011110001: out = 32'b00000000000000000111100100001111;
            12'b000011110010: out = 32'b00000000000000000111100110010000;
            12'b000011110011: out = 32'b00000000000000000111101000010010;
            12'b000011110100: out = 32'b00000000000000000111101010010100;
            12'b000011110101: out = 32'b00000000000000000111101100010110;
            12'b000011110110: out = 32'b00000000000000000111101110011000;
            12'b000011110111: out = 32'b00000000000000000111110000011010;
            12'b000011111000: out = 32'b00000000000000000111110010011100;
            12'b000011111001: out = 32'b00000000000000000111110100011101;
            12'b000011111010: out = 32'b00000000000000000111110110011111;
            12'b000011111011: out = 32'b00000000000000000111111000100001;
            12'b000011111100: out = 32'b00000000000000000111111010100011;
            12'b000011111101: out = 32'b00000000000000000111111100100101;
            12'b000011111110: out = 32'b00000000000000000111111110100111;
            12'b000011111111: out = 32'b00000000000000001000000000101001;
            12'b000100000000: out = 32'b00000000000000001000000010101011;
            12'b000100000001: out = 32'b00000000000000001000000100101101;
            12'b000100000010: out = 32'b00000000000000001000000110101111;
            12'b000100000011: out = 32'b00000000000000001000001000110001;
            12'b000100000100: out = 32'b00000000000000001000001010110011;
            12'b000100000101: out = 32'b00000000000000001000001100110110;
            12'b000100000110: out = 32'b00000000000000001000001110111000;
            12'b000100000111: out = 32'b00000000000000001000010000111010;
            12'b000100001000: out = 32'b00000000000000001000010010111100;
            12'b000100001001: out = 32'b00000000000000001000010100111110;
            12'b000100001010: out = 32'b00000000000000001000010111000000;
            12'b000100001011: out = 32'b00000000000000001000011001000010;
            12'b000100001100: out = 32'b00000000000000001000011011000101;
            12'b000100001101: out = 32'b00000000000000001000011101000111;
            12'b000100001110: out = 32'b00000000000000001000011111001001;
            12'b000100001111: out = 32'b00000000000000001000100001001011;
            12'b000100010000: out = 32'b00000000000000001000100011001110;
            12'b000100010001: out = 32'b00000000000000001000100101010000;
            12'b000100010010: out = 32'b00000000000000001000100111010010;
            12'b000100010011: out = 32'b00000000000000001000101001010101;
            12'b000100010100: out = 32'b00000000000000001000101011010111;
            12'b000100010101: out = 32'b00000000000000001000101101011001;
            12'b000100010110: out = 32'b00000000000000001000101111011100;
            12'b000100010111: out = 32'b00000000000000001000110001011110;
            12'b000100011000: out = 32'b00000000000000001000110011100000;
            12'b000100011001: out = 32'b00000000000000001000110101100011;
            12'b000100011010: out = 32'b00000000000000001000110111100101;
            12'b000100011011: out = 32'b00000000000000001000111001101000;
            12'b000100011100: out = 32'b00000000000000001000111011101010;
            12'b000100011101: out = 32'b00000000000000001000111101101101;
            12'b000100011110: out = 32'b00000000000000001000111111101111;
            12'b000100011111: out = 32'b00000000000000001001000001110010;
            12'b000100100000: out = 32'b00000000000000001001000011110100;
            12'b000100100001: out = 32'b00000000000000001001000101110111;
            12'b000100100010: out = 32'b00000000000000001001000111111010;
            12'b000100100011: out = 32'b00000000000000001001001001111100;
            12'b000100100100: out = 32'b00000000000000001001001011111111;
            12'b000100100101: out = 32'b00000000000000001001001110000001;
            12'b000100100110: out = 32'b00000000000000001001010000000100;
            12'b000100100111: out = 32'b00000000000000001001010010000111;
            12'b000100101000: out = 32'b00000000000000001001010100001010;
            12'b000100101001: out = 32'b00000000000000001001010110001100;
            12'b000100101010: out = 32'b00000000000000001001011000001111;
            12'b000100101011: out = 32'b00000000000000001001011010010010;
            12'b000100101100: out = 32'b00000000000000001001011100010101;
            12'b000100101101: out = 32'b00000000000000001001011110010111;
            12'b000100101110: out = 32'b00000000000000001001100000011010;
            12'b000100101111: out = 32'b00000000000000001001100010011101;
            12'b000100110000: out = 32'b00000000000000001001100100100000;
            12'b000100110001: out = 32'b00000000000000001001100110100011;
            12'b000100110010: out = 32'b00000000000000001001101000100110;
            12'b000100110011: out = 32'b00000000000000001001101010101001;
            12'b000100110100: out = 32'b00000000000000001001101100101011;
            12'b000100110101: out = 32'b00000000000000001001101110101110;
            12'b000100110110: out = 32'b00000000000000001001110000110001;
            12'b000100110111: out = 32'b00000000000000001001110010110100;
            12'b000100111000: out = 32'b00000000000000001001110100110111;
            12'b000100111001: out = 32'b00000000000000001001110110111010;
            12'b000100111010: out = 32'b00000000000000001001111000111101;
            12'b000100111011: out = 32'b00000000000000001001111011000000;
            12'b000100111100: out = 32'b00000000000000001001111101000100;
            12'b000100111101: out = 32'b00000000000000001001111111000111;
            12'b000100111110: out = 32'b00000000000000001010000001001010;
            12'b000100111111: out = 32'b00000000000000001010000011001101;
            12'b000101000000: out = 32'b00000000000000001010000101010000;
            12'b000101000001: out = 32'b00000000000000001010000111010011;
            12'b000101000010: out = 32'b00000000000000001010001001010111;
            12'b000101000011: out = 32'b00000000000000001010001011011010;
            12'b000101000100: out = 32'b00000000000000001010001101011101;
            12'b000101000101: out = 32'b00000000000000001010001111100000;
            12'b000101000110: out = 32'b00000000000000001010010001100100;
            12'b000101000111: out = 32'b00000000000000001010010011100111;
            12'b000101001000: out = 32'b00000000000000001010010101101010;
            12'b000101001001: out = 32'b00000000000000001010010111101110;
            12'b000101001010: out = 32'b00000000000000001010011001110001;
            12'b000101001011: out = 32'b00000000000000001010011011110100;
            12'b000101001100: out = 32'b00000000000000001010011101111000;
            12'b000101001101: out = 32'b00000000000000001010011111111011;
            12'b000101001110: out = 32'b00000000000000001010100001111111;
            12'b000101001111: out = 32'b00000000000000001010100100000010;
            12'b000101010000: out = 32'b00000000000000001010100110000110;
            12'b000101010001: out = 32'b00000000000000001010101000001001;
            12'b000101010010: out = 32'b00000000000000001010101010001101;
            12'b000101010011: out = 32'b00000000000000001010101100010000;
            12'b000101010100: out = 32'b00000000000000001010101110010100;
            12'b000101010101: out = 32'b00000000000000001010110000010111;
            12'b000101010110: out = 32'b00000000000000001010110010011011;
            12'b000101010111: out = 32'b00000000000000001010110100011111;
            12'b000101011000: out = 32'b00000000000000001010110110100010;
            12'b000101011001: out = 32'b00000000000000001010111000100110;
            12'b000101011010: out = 32'b00000000000000001010111010101010;
            12'b000101011011: out = 32'b00000000000000001010111100101101;
            12'b000101011100: out = 32'b00000000000000001010111110110001;
            12'b000101011101: out = 32'b00000000000000001011000000110101;
            12'b000101011110: out = 32'b00000000000000001011000010111001;
            12'b000101011111: out = 32'b00000000000000001011000100111101;
            12'b000101100000: out = 32'b00000000000000001011000111000000;
            12'b000101100001: out = 32'b00000000000000001011001001000100;
            12'b000101100010: out = 32'b00000000000000001011001011001000;
            12'b000101100011: out = 32'b00000000000000001011001101001100;
            12'b000101100100: out = 32'b00000000000000001011001111010000;
            12'b000101100101: out = 32'b00000000000000001011010001010100;
            12'b000101100110: out = 32'b00000000000000001011010011011000;
            12'b000101100111: out = 32'b00000000000000001011010101011100;
            12'b000101101000: out = 32'b00000000000000001011010111100000;
            12'b000101101001: out = 32'b00000000000000001011011001100100;
            12'b000101101010: out = 32'b00000000000000001011011011101000;
            12'b000101101011: out = 32'b00000000000000001011011101101100;
            12'b000101101100: out = 32'b00000000000000001011011111110000;
            12'b000101101101: out = 32'b00000000000000001011100001110101;
            12'b000101101110: out = 32'b00000000000000001011100011111001;
            12'b000101101111: out = 32'b00000000000000001011100101111101;
            12'b000101110000: out = 32'b00000000000000001011101000000001;
            12'b000101110001: out = 32'b00000000000000001011101010000101;
            12'b000101110010: out = 32'b00000000000000001011101100001010;
            12'b000101110011: out = 32'b00000000000000001011101110001110;
            12'b000101110100: out = 32'b00000000000000001011110000010010;
            12'b000101110101: out = 32'b00000000000000001011110010010111;
            12'b000101110110: out = 32'b00000000000000001011110100011011;
            12'b000101110111: out = 32'b00000000000000001011110110011111;
            12'b000101111000: out = 32'b00000000000000001011111000100100;
            12'b000101111001: out = 32'b00000000000000001011111010101000;
            12'b000101111010: out = 32'b00000000000000001011111100101101;
            12'b000101111011: out = 32'b00000000000000001011111110110001;
            12'b000101111100: out = 32'b00000000000000001100000000110101;
            12'b000101111101: out = 32'b00000000000000001100000010111010;
            12'b000101111110: out = 32'b00000000000000001100000100111111;
            12'b000101111111: out = 32'b00000000000000001100000111000011;
            12'b000110000000: out = 32'b00000000000000001100001001001000;
            12'b000110000001: out = 32'b00000000000000001100001011001100;
            12'b000110000010: out = 32'b00000000000000001100001101010001;
            12'b000110000011: out = 32'b00000000000000001100001111010110;
            12'b000110000100: out = 32'b00000000000000001100010001011010;
            12'b000110000101: out = 32'b00000000000000001100010011011111;
            12'b000110000110: out = 32'b00000000000000001100010101100100;
            12'b000110000111: out = 32'b00000000000000001100010111101001;
            12'b000110001000: out = 32'b00000000000000001100011001101101;
            12'b000110001001: out = 32'b00000000000000001100011011110010;
            12'b000110001010: out = 32'b00000000000000001100011101110111;
            12'b000110001011: out = 32'b00000000000000001100011111111100;
            12'b000110001100: out = 32'b00000000000000001100100010000001;
            12'b000110001101: out = 32'b00000000000000001100100100000110;
            12'b000110001110: out = 32'b00000000000000001100100110001011;
            12'b000110001111: out = 32'b00000000000000001100101000010000;
            12'b000110010000: out = 32'b00000000000000001100101010010101;
            12'b000110010001: out = 32'b00000000000000001100101100011010;
            12'b000110010010: out = 32'b00000000000000001100101110011111;
            12'b000110010011: out = 32'b00000000000000001100110000100100;
            12'b000110010100: out = 32'b00000000000000001100110010101001;
            12'b000110010101: out = 32'b00000000000000001100110100101110;
            12'b000110010110: out = 32'b00000000000000001100110110110011;
            12'b000110010111: out = 32'b00000000000000001100111000111000;
            12'b000110011000: out = 32'b00000000000000001100111010111110;
            12'b000110011001: out = 32'b00000000000000001100111101000011;
            12'b000110011010: out = 32'b00000000000000001100111111001000;
            12'b000110011011: out = 32'b00000000000000001101000001001101;
            12'b000110011100: out = 32'b00000000000000001101000011010011;
            12'b000110011101: out = 32'b00000000000000001101000101011000;
            12'b000110011110: out = 32'b00000000000000001101000111011101;
            12'b000110011111: out = 32'b00000000000000001101001001100011;
            12'b000110100000: out = 32'b00000000000000001101001011101000;
            12'b000110100001: out = 32'b00000000000000001101001101101110;
            12'b000110100010: out = 32'b00000000000000001101001111110011;
            12'b000110100011: out = 32'b00000000000000001101010001111001;
            12'b000110100100: out = 32'b00000000000000001101010011111110;
            12'b000110100101: out = 32'b00000000000000001101010110000100;
            12'b000110100110: out = 32'b00000000000000001101011000001001;
            12'b000110100111: out = 32'b00000000000000001101011010001111;
            12'b000110101000: out = 32'b00000000000000001101011100010100;
            12'b000110101001: out = 32'b00000000000000001101011110011010;
            12'b000110101010: out = 32'b00000000000000001101100000100000;
            12'b000110101011: out = 32'b00000000000000001101100010100101;
            12'b000110101100: out = 32'b00000000000000001101100100101011;
            12'b000110101101: out = 32'b00000000000000001101100110110001;
            12'b000110101110: out = 32'b00000000000000001101101000110111;
            12'b000110101111: out = 32'b00000000000000001101101010111101;
            12'b000110110000: out = 32'b00000000000000001101101101000010;
            12'b000110110001: out = 32'b00000000000000001101101111001000;
            12'b000110110010: out = 32'b00000000000000001101110001001110;
            12'b000110110011: out = 32'b00000000000000001101110011010100;
            12'b000110110100: out = 32'b00000000000000001101110101011010;
            12'b000110110101: out = 32'b00000000000000001101110111100000;
            12'b000110110110: out = 32'b00000000000000001101111001100110;
            12'b000110110111: out = 32'b00000000000000001101111011101100;
            12'b000110111000: out = 32'b00000000000000001101111101110010;
            12'b000110111001: out = 32'b00000000000000001101111111111000;
            12'b000110111010: out = 32'b00000000000000001110000001111111;
            12'b000110111011: out = 32'b00000000000000001110000100000101;
            12'b000110111100: out = 32'b00000000000000001110000110001011;
            12'b000110111101: out = 32'b00000000000000001110001000010001;
            12'b000110111110: out = 32'b00000000000000001110001010010111;
            12'b000110111111: out = 32'b00000000000000001110001100011110;
            12'b000111000000: out = 32'b00000000000000001110001110100100;
            12'b000111000001: out = 32'b00000000000000001110010000101010;
            12'b000111000010: out = 32'b00000000000000001110010010110001;
            12'b000111000011: out = 32'b00000000000000001110010100110111;
            12'b000111000100: out = 32'b00000000000000001110010110111110;
            12'b000111000101: out = 32'b00000000000000001110011001000100;
            12'b000111000110: out = 32'b00000000000000001110011011001011;
            12'b000111000111: out = 32'b00000000000000001110011101010001;
            12'b000111001000: out = 32'b00000000000000001110011111011000;
            12'b000111001001: out = 32'b00000000000000001110100001011110;
            12'b000111001010: out = 32'b00000000000000001110100011100101;
            12'b000111001011: out = 32'b00000000000000001110100101101011;
            12'b000111001100: out = 32'b00000000000000001110100111110010;
            12'b000111001101: out = 32'b00000000000000001110101001111001;
            12'b000111001110: out = 32'b00000000000000001110101011111111;
            12'b000111001111: out = 32'b00000000000000001110101110000110;
            12'b000111010000: out = 32'b00000000000000001110110000001101;
            12'b000111010001: out = 32'b00000000000000001110110010010100;
            12'b000111010010: out = 32'b00000000000000001110110100011011;
            12'b000111010011: out = 32'b00000000000000001110110110100010;
            12'b000111010100: out = 32'b00000000000000001110111000101000;
            12'b000111010101: out = 32'b00000000000000001110111010101111;
            12'b000111010110: out = 32'b00000000000000001110111100110110;
            12'b000111010111: out = 32'b00000000000000001110111110111101;
            12'b000111011000: out = 32'b00000000000000001111000001000100;
            12'b000111011001: out = 32'b00000000000000001111000011001011;
            12'b000111011010: out = 32'b00000000000000001111000101010011;
            12'b000111011011: out = 32'b00000000000000001111000111011010;
            12'b000111011100: out = 32'b00000000000000001111001001100001;
            12'b000111011101: out = 32'b00000000000000001111001011101000;
            12'b000111011110: out = 32'b00000000000000001111001101101111;
            12'b000111011111: out = 32'b00000000000000001111001111110111;
            12'b000111100000: out = 32'b00000000000000001111010001111110;
            12'b000111100001: out = 32'b00000000000000001111010100000101;
            12'b000111100010: out = 32'b00000000000000001111010110001100;
            12'b000111100011: out = 32'b00000000000000001111011000010100;
            12'b000111100100: out = 32'b00000000000000001111011010011011;
            12'b000111100101: out = 32'b00000000000000001111011100100011;
            12'b000111100110: out = 32'b00000000000000001111011110101010;
            12'b000111100111: out = 32'b00000000000000001111100000110010;
            12'b000111101000: out = 32'b00000000000000001111100010111001;
            12'b000111101001: out = 32'b00000000000000001111100101000001;
            12'b000111101010: out = 32'b00000000000000001111100111001000;
            12'b000111101011: out = 32'b00000000000000001111101001010000;
            12'b000111101100: out = 32'b00000000000000001111101011011000;
            12'b000111101101: out = 32'b00000000000000001111101101011111;
            12'b000111101110: out = 32'b00000000000000001111101111100111;
            12'b000111101111: out = 32'b00000000000000001111110001101111;
            12'b000111110000: out = 32'b00000000000000001111110011110111;
            12'b000111110001: out = 32'b00000000000000001111110101111110;
            12'b000111110010: out = 32'b00000000000000001111111000000110;
            12'b000111110011: out = 32'b00000000000000001111111010001110;
            12'b000111110100: out = 32'b00000000000000001111111100010110;
            12'b000111110101: out = 32'b00000000000000001111111110011110;
            12'b000111110110: out = 32'b00000000000000010000000000100110;
            12'b000111110111: out = 32'b00000000000000010000000010101110;
            12'b000111111000: out = 32'b00000000000000010000000100110110;
            12'b000111111001: out = 32'b00000000000000010000000110111110;
            12'b000111111010: out = 32'b00000000000000010000001001000110;
            12'b000111111011: out = 32'b00000000000000010000001011001111;
            12'b000111111100: out = 32'b00000000000000010000001101010111;
            12'b000111111101: out = 32'b00000000000000010000001111011111;
            12'b000111111110: out = 32'b00000000000000010000010001100111;
            12'b000111111111: out = 32'b00000000000000010000010011110000;
            12'b001000000000: out = 32'b00000000000000010000010101111000;
            12'b001000000001: out = 32'b00000000000000010000011000000000;
            12'b001000000010: out = 32'b00000000000000010000011010001001;
            12'b001000000011: out = 32'b00000000000000010000011100010001;
            12'b001000000100: out = 32'b00000000000000010000011110011010;
            12'b001000000101: out = 32'b00000000000000010000100000100010;
            12'b001000000110: out = 32'b00000000000000010000100010101011;
            12'b001000000111: out = 32'b00000000000000010000100100110011;
            12'b001000001000: out = 32'b00000000000000010000100110111100;
            12'b001000001001: out = 32'b00000000000000010000101001000100;
            12'b001000001010: out = 32'b00000000000000010000101011001101;
            12'b001000001011: out = 32'b00000000000000010000101101010110;
            12'b001000001100: out = 32'b00000000000000010000101111011110;
            12'b001000001101: out = 32'b00000000000000010000110001100111;
            12'b001000001110: out = 32'b00000000000000010000110011110000;
            12'b001000001111: out = 32'b00000000000000010000110101111001;
            12'b001000010000: out = 32'b00000000000000010000111000000010;
            12'b001000010001: out = 32'b00000000000000010000111010001011;
            12'b001000010010: out = 32'b00000000000000010000111100010100;
            12'b001000010011: out = 32'b00000000000000010000111110011101;
            12'b001000010100: out = 32'b00000000000000010001000000100110;
            12'b001000010101: out = 32'b00000000000000010001000010101111;
            12'b001000010110: out = 32'b00000000000000010001000100111000;
            12'b001000010111: out = 32'b00000000000000010001000111000001;
            12'b001000011000: out = 32'b00000000000000010001001001001010;
            12'b001000011001: out = 32'b00000000000000010001001011010011;
            12'b001000011010: out = 32'b00000000000000010001001101011101;
            12'b001000011011: out = 32'b00000000000000010001001111100110;
            12'b001000011100: out = 32'b00000000000000010001010001101111;
            12'b001000011101: out = 32'b00000000000000010001010011111000;
            12'b001000011110: out = 32'b00000000000000010001010110000010;
            12'b001000011111: out = 32'b00000000000000010001011000001011;
            12'b001000100000: out = 32'b00000000000000010001011010010101;
            12'b001000100001: out = 32'b00000000000000010001011100011110;
            12'b001000100010: out = 32'b00000000000000010001011110101000;
            12'b001000100011: out = 32'b00000000000000010001100000110001;
            12'b001000100100: out = 32'b00000000000000010001100010111011;
            12'b001000100101: out = 32'b00000000000000010001100101000101;
            12'b001000100110: out = 32'b00000000000000010001100111001110;
            12'b001000100111: out = 32'b00000000000000010001101001011000;
            12'b001000101000: out = 32'b00000000000000010001101011100010;
            12'b001000101001: out = 32'b00000000000000010001101101101011;
            12'b001000101010: out = 32'b00000000000000010001101111110101;
            12'b001000101011: out = 32'b00000000000000010001110001111111;
            12'b001000101100: out = 32'b00000000000000010001110100001001;
            12'b001000101101: out = 32'b00000000000000010001110110010011;
            12'b001000101110: out = 32'b00000000000000010001111000011101;
            12'b001000101111: out = 32'b00000000000000010001111010100111;
            12'b001000110000: out = 32'b00000000000000010001111100110001;
            12'b001000110001: out = 32'b00000000000000010001111110111011;
            12'b001000110010: out = 32'b00000000000000010010000001000101;
            12'b001000110011: out = 32'b00000000000000010010000011001111;
            12'b001000110100: out = 32'b00000000000000010010000101011010;
            12'b001000110101: out = 32'b00000000000000010010000111100100;
            12'b001000110110: out = 32'b00000000000000010010001001101110;
            12'b001000110111: out = 32'b00000000000000010010001011111000;
            12'b001000111000: out = 32'b00000000000000010010001110000011;
            12'b001000111001: out = 32'b00000000000000010010010000001101;
            12'b001000111010: out = 32'b00000000000000010010010010011000;
            12'b001000111011: out = 32'b00000000000000010010010100100010;
            12'b001000111100: out = 32'b00000000000000010010010110101101;
            12'b001000111101: out = 32'b00000000000000010010011000110111;
            12'b001000111110: out = 32'b00000000000000010010011011000010;
            12'b001000111111: out = 32'b00000000000000010010011101001100;
            12'b001001000000: out = 32'b00000000000000010010011111010111;
            12'b001001000001: out = 32'b00000000000000010010100001100010;
            12'b001001000010: out = 32'b00000000000000010010100011101100;
            12'b001001000011: out = 32'b00000000000000010010100101110111;
            12'b001001000100: out = 32'b00000000000000010010101000000010;
            12'b001001000101: out = 32'b00000000000000010010101010001101;
            12'b001001000110: out = 32'b00000000000000010010101100011000;
            12'b001001000111: out = 32'b00000000000000010010101110100011;
            12'b001001001000: out = 32'b00000000000000010010110000101110;
            12'b001001001001: out = 32'b00000000000000010010110010111001;
            12'b001001001010: out = 32'b00000000000000010010110101000100;
            12'b001001001011: out = 32'b00000000000000010010110111001111;
            12'b001001001100: out = 32'b00000000000000010010111001011010;
            12'b001001001101: out = 32'b00000000000000010010111011100101;
            12'b001001001110: out = 32'b00000000000000010010111101110000;
            12'b001001001111: out = 32'b00000000000000010010111111111100;
            12'b001001010000: out = 32'b00000000000000010011000010000111;
            12'b001001010001: out = 32'b00000000000000010011000100010010;
            12'b001001010010: out = 32'b00000000000000010011000110011110;
            12'b001001010011: out = 32'b00000000000000010011001000101001;
            12'b001001010100: out = 32'b00000000000000010011001010110101;
            12'b001001010101: out = 32'b00000000000000010011001101000000;
            12'b001001010110: out = 32'b00000000000000010011001111001100;
            12'b001001010111: out = 32'b00000000000000010011010001010111;
            12'b001001011000: out = 32'b00000000000000010011010011100011;
            12'b001001011001: out = 32'b00000000000000010011010101101111;
            12'b001001011010: out = 32'b00000000000000010011010111111010;
            12'b001001011011: out = 32'b00000000000000010011011010000110;
            12'b001001011100: out = 32'b00000000000000010011011100010010;
            12'b001001011101: out = 32'b00000000000000010011011110011110;
            12'b001001011110: out = 32'b00000000000000010011100000101010;
            12'b001001011111: out = 32'b00000000000000010011100010110101;
            12'b001001100000: out = 32'b00000000000000010011100101000001;
            12'b001001100001: out = 32'b00000000000000010011100111001101;
            12'b001001100010: out = 32'b00000000000000010011101001011001;
            12'b001001100011: out = 32'b00000000000000010011101011100110;
            12'b001001100100: out = 32'b00000000000000010011101101110010;
            12'b001001100101: out = 32'b00000000000000010011101111111110;
            12'b001001100110: out = 32'b00000000000000010011110010001010;
            12'b001001100111: out = 32'b00000000000000010011110100010110;
            12'b001001101000: out = 32'b00000000000000010011110110100011;
            12'b001001101001: out = 32'b00000000000000010011111000101111;
            12'b001001101010: out = 32'b00000000000000010011111010111011;
            12'b001001101011: out = 32'b00000000000000010011111101001000;
            12'b001001101100: out = 32'b00000000000000010011111111010100;
            12'b001001101101: out = 32'b00000000000000010100000001100001;
            12'b001001101110: out = 32'b00000000000000010100000011101101;
            12'b001001101111: out = 32'b00000000000000010100000101111010;
            12'b001001110000: out = 32'b00000000000000010100001000000110;
            12'b001001110001: out = 32'b00000000000000010100001010010011;
            12'b001001110010: out = 32'b00000000000000010100001100100000;
            12'b001001110011: out = 32'b00000000000000010100001110101101;
            12'b001001110100: out = 32'b00000000000000010100010000111001;
            12'b001001110101: out = 32'b00000000000000010100010011000110;
            12'b001001110110: out = 32'b00000000000000010100010101010011;
            12'b001001110111: out = 32'b00000000000000010100010111100000;
            12'b001001111000: out = 32'b00000000000000010100011001101101;
            12'b001001111001: out = 32'b00000000000000010100011011111010;
            12'b001001111010: out = 32'b00000000000000010100011110000111;
            12'b001001111011: out = 32'b00000000000000010100100000010100;
            12'b001001111100: out = 32'b00000000000000010100100010100010;
            12'b001001111101: out = 32'b00000000000000010100100100101111;
            12'b001001111110: out = 32'b00000000000000010100100110111100;
            12'b001001111111: out = 32'b00000000000000010100101001001001;
            12'b001010000000: out = 32'b00000000000000010100101011010111;
            12'b001010000001: out = 32'b00000000000000010100101101100100;
            12'b001010000010: out = 32'b00000000000000010100101111110001;
            12'b001010000011: out = 32'b00000000000000010100110001111111;
            12'b001010000100: out = 32'b00000000000000010100110100001100;
            12'b001010000101: out = 32'b00000000000000010100110110011010;
            12'b001010000110: out = 32'b00000000000000010100111000101000;
            12'b001010000111: out = 32'b00000000000000010100111010110101;
            12'b001010001000: out = 32'b00000000000000010100111101000011;
            12'b001010001001: out = 32'b00000000000000010100111111010001;
            12'b001010001010: out = 32'b00000000000000010101000001011110;
            12'b001010001011: out = 32'b00000000000000010101000011101100;
            12'b001010001100: out = 32'b00000000000000010101000101111010;
            12'b001010001101: out = 32'b00000000000000010101001000001000;
            12'b001010001110: out = 32'b00000000000000010101001010010110;
            12'b001010001111: out = 32'b00000000000000010101001100100100;
            12'b001010010000: out = 32'b00000000000000010101001110110010;
            12'b001010010001: out = 32'b00000000000000010101010001000000;
            12'b001010010010: out = 32'b00000000000000010101010011001110;
            12'b001010010011: out = 32'b00000000000000010101010101011101;
            12'b001010010100: out = 32'b00000000000000010101010111101011;
            12'b001010010101: out = 32'b00000000000000010101011001111001;
            12'b001010010110: out = 32'b00000000000000010101011100001000;
            12'b001010010111: out = 32'b00000000000000010101011110010110;
            12'b001010011000: out = 32'b00000000000000010101100000100100;
            12'b001010011001: out = 32'b00000000000000010101100010110011;
            12'b001010011010: out = 32'b00000000000000010101100101000001;
            12'b001010011011: out = 32'b00000000000000010101100111010000;
            12'b001010011100: out = 32'b00000000000000010101101001011111;
            12'b001010011101: out = 32'b00000000000000010101101011101101;
            12'b001010011110: out = 32'b00000000000000010101101101111100;
            12'b001010011111: out = 32'b00000000000000010101110000001011;
            12'b001010100000: out = 32'b00000000000000010101110010011010;
            12'b001010100001: out = 32'b00000000000000010101110100101000;
            12'b001010100010: out = 32'b00000000000000010101110110110111;
            12'b001010100011: out = 32'b00000000000000010101111001000110;
            12'b001010100100: out = 32'b00000000000000010101111011010101;
            12'b001010100101: out = 32'b00000000000000010101111101100100;
            12'b001010100110: out = 32'b00000000000000010101111111110011;
            12'b001010100111: out = 32'b00000000000000010110000010000011;
            12'b001010101000: out = 32'b00000000000000010110000100010010;
            12'b001010101001: out = 32'b00000000000000010110000110100001;
            12'b001010101010: out = 32'b00000000000000010110001000110000;
            12'b001010101011: out = 32'b00000000000000010110001011000000;
            12'b001010101100: out = 32'b00000000000000010110001101001111;
            12'b001010101101: out = 32'b00000000000000010110001111011110;
            12'b001010101110: out = 32'b00000000000000010110010001101110;
            12'b001010101111: out = 32'b00000000000000010110010011111101;
            12'b001010110000: out = 32'b00000000000000010110010110001101;
            12'b001010110001: out = 32'b00000000000000010110011000011101;
            12'b001010110010: out = 32'b00000000000000010110011010101100;
            12'b001010110011: out = 32'b00000000000000010110011100111100;
            12'b001010110100: out = 32'b00000000000000010110011111001100;
            12'b001010110101: out = 32'b00000000000000010110100001011100;
            12'b001010110110: out = 32'b00000000000000010110100011101100;
            12'b001010110111: out = 32'b00000000000000010110100101111011;
            12'b001010111000: out = 32'b00000000000000010110101000001011;
            12'b001010111001: out = 32'b00000000000000010110101010011011;
            12'b001010111010: out = 32'b00000000000000010110101100101100;
            12'b001010111011: out = 32'b00000000000000010110101110111100;
            12'b001010111100: out = 32'b00000000000000010110110001001100;
            12'b001010111101: out = 32'b00000000000000010110110011011100;
            12'b001010111110: out = 32'b00000000000000010110110101101100;
            12'b001010111111: out = 32'b00000000000000010110110111111101;
            12'b001011000000: out = 32'b00000000000000010110111010001101;
            12'b001011000001: out = 32'b00000000000000010110111100011101;
            12'b001011000010: out = 32'b00000000000000010110111110101110;
            12'b001011000011: out = 32'b00000000000000010111000000111110;
            12'b001011000100: out = 32'b00000000000000010111000011001111;
            12'b001011000101: out = 32'b00000000000000010111000101100000;
            12'b001011000110: out = 32'b00000000000000010111000111110000;
            12'b001011000111: out = 32'b00000000000000010111001010000001;
            12'b001011001000: out = 32'b00000000000000010111001100010010;
            12'b001011001001: out = 32'b00000000000000010111001110100011;
            12'b001011001010: out = 32'b00000000000000010111010000110100;
            12'b001011001011: out = 32'b00000000000000010111010011000101;
            12'b001011001100: out = 32'b00000000000000010111010101010110;
            12'b001011001101: out = 32'b00000000000000010111010111100111;
            12'b001011001110: out = 32'b00000000000000010111011001111000;
            12'b001011001111: out = 32'b00000000000000010111011100001001;
            12'b001011010000: out = 32'b00000000000000010111011110011010;
            12'b001011010001: out = 32'b00000000000000010111100000101011;
            12'b001011010010: out = 32'b00000000000000010111100010111101;
            12'b001011010011: out = 32'b00000000000000010111100101001110;
            12'b001011010100: out = 32'b00000000000000010111100111011111;
            12'b001011010101: out = 32'b00000000000000010111101001110001;
            12'b001011010110: out = 32'b00000000000000010111101100000010;
            12'b001011010111: out = 32'b00000000000000010111101110010100;
            12'b001011011000: out = 32'b00000000000000010111110000100101;
            12'b001011011001: out = 32'b00000000000000010111110010110111;
            12'b001011011010: out = 32'b00000000000000010111110101001001;
            12'b001011011011: out = 32'b00000000000000010111110111011011;
            12'b001011011100: out = 32'b00000000000000010111111001101100;
            12'b001011011101: out = 32'b00000000000000010111111011111110;
            12'b001011011110: out = 32'b00000000000000010111111110010000;
            12'b001011011111: out = 32'b00000000000000011000000000100010;
            12'b001011100000: out = 32'b00000000000000011000000010110100;
            12'b001011100001: out = 32'b00000000000000011000000101000110;
            12'b001011100010: out = 32'b00000000000000011000000111011000;
            12'b001011100011: out = 32'b00000000000000011000001001101011;
            12'b001011100100: out = 32'b00000000000000011000001011111101;
            12'b001011100101: out = 32'b00000000000000011000001110001111;
            12'b001011100110: out = 32'b00000000000000011000010000100010;
            12'b001011100111: out = 32'b00000000000000011000010010110100;
            12'b001011101000: out = 32'b00000000000000011000010101000110;
            12'b001011101001: out = 32'b00000000000000011000010111011001;
            12'b001011101010: out = 32'b00000000000000011000011001101100;
            12'b001011101011: out = 32'b00000000000000011000011011111110;
            12'b001011101100: out = 32'b00000000000000011000011110010001;
            12'b001011101101: out = 32'b00000000000000011000100000100100;
            12'b001011101110: out = 32'b00000000000000011000100010110110;
            12'b001011101111: out = 32'b00000000000000011000100101001001;
            12'b001011110000: out = 32'b00000000000000011000100111011100;
            12'b001011110001: out = 32'b00000000000000011000101001101111;
            12'b001011110010: out = 32'b00000000000000011000101100000010;
            12'b001011110011: out = 32'b00000000000000011000101110010101;
            12'b001011110100: out = 32'b00000000000000011000110000101000;
            12'b001011110101: out = 32'b00000000000000011000110010111100;
            12'b001011110110: out = 32'b00000000000000011000110101001111;
            12'b001011110111: out = 32'b00000000000000011000110111100010;
            12'b001011111000: out = 32'b00000000000000011000111001110101;
            12'b001011111001: out = 32'b00000000000000011000111100001001;
            12'b001011111010: out = 32'b00000000000000011000111110011100;
            12'b001011111011: out = 32'b00000000000000011001000000110000;
            12'b001011111100: out = 32'b00000000000000011001000011000011;
            12'b001011111101: out = 32'b00000000000000011001000101010111;
            12'b001011111110: out = 32'b00000000000000011001000111101011;
            12'b001011111111: out = 32'b00000000000000011001001001111111;
            12'b001100000000: out = 32'b00000000000000011001001100010010;
            12'b001100000001: out = 32'b00000000000000011001001110100110;
            12'b001100000010: out = 32'b00000000000000011001010000111010;
            12'b001100000011: out = 32'b00000000000000011001010011001110;
            12'b001100000100: out = 32'b00000000000000011001010101100010;
            12'b001100000101: out = 32'b00000000000000011001010111110110;
            12'b001100000110: out = 32'b00000000000000011001011010001010;
            12'b001100000111: out = 32'b00000000000000011001011100011111;
            12'b001100001000: out = 32'b00000000000000011001011110110011;
            12'b001100001001: out = 32'b00000000000000011001100001000111;
            12'b001100001010: out = 32'b00000000000000011001100011011100;
            12'b001100001011: out = 32'b00000000000000011001100101110000;
            12'b001100001100: out = 32'b00000000000000011001101000000100;
            12'b001100001101: out = 32'b00000000000000011001101010011001;
            12'b001100001110: out = 32'b00000000000000011001101100101110;
            12'b001100001111: out = 32'b00000000000000011001101111000010;
            12'b001100010000: out = 32'b00000000000000011001110001010111;
            12'b001100010001: out = 32'b00000000000000011001110011101100;
            12'b001100010010: out = 32'b00000000000000011001110110000001;
            12'b001100010011: out = 32'b00000000000000011001111000010110;
            12'b001100010100: out = 32'b00000000000000011001111010101011;
            12'b001100010101: out = 32'b00000000000000011001111101000000;
            12'b001100010110: out = 32'b00000000000000011001111111010101;
            12'b001100010111: out = 32'b00000000000000011010000001101010;
            12'b001100011000: out = 32'b00000000000000011010000011111111;
            12'b001100011001: out = 32'b00000000000000011010000110010100;
            12'b001100011010: out = 32'b00000000000000011010001000101010;
            12'b001100011011: out = 32'b00000000000000011010001010111111;
            12'b001100011100: out = 32'b00000000000000011010001101010100;
            12'b001100011101: out = 32'b00000000000000011010001111101010;
            12'b001100011110: out = 32'b00000000000000011010010001111111;
            12'b001100011111: out = 32'b00000000000000011010010100010101;
            12'b001100100000: out = 32'b00000000000000011010010110101011;
            12'b001100100001: out = 32'b00000000000000011010011001000000;
            12'b001100100010: out = 32'b00000000000000011010011011010110;
            12'b001100100011: out = 32'b00000000000000011010011101101100;
            12'b001100100100: out = 32'b00000000000000011010100000000010;
            12'b001100100101: out = 32'b00000000000000011010100010011000;
            12'b001100100110: out = 32'b00000000000000011010100100101110;
            12'b001100100111: out = 32'b00000000000000011010100111000100;
            12'b001100101000: out = 32'b00000000000000011010101001011010;
            12'b001100101001: out = 32'b00000000000000011010101011110000;
            12'b001100101010: out = 32'b00000000000000011010101110000111;
            12'b001100101011: out = 32'b00000000000000011010110000011101;
            12'b001100101100: out = 32'b00000000000000011010110010110011;
            12'b001100101101: out = 32'b00000000000000011010110101001010;
            12'b001100101110: out = 32'b00000000000000011010110111100000;
            12'b001100101111: out = 32'b00000000000000011010111001110111;
            12'b001100110000: out = 32'b00000000000000011010111100001110;
            12'b001100110001: out = 32'b00000000000000011010111110100100;
            12'b001100110010: out = 32'b00000000000000011011000000111011;
            12'b001100110011: out = 32'b00000000000000011011000011010010;
            12'b001100110100: out = 32'b00000000000000011011000101101001;
            12'b001100110101: out = 32'b00000000000000011011001000000000;
            12'b001100110110: out = 32'b00000000000000011011001010010111;
            12'b001100110111: out = 32'b00000000000000011011001100101110;
            12'b001100111000: out = 32'b00000000000000011011001111000101;
            12'b001100111001: out = 32'b00000000000000011011010001011100;
            12'b001100111010: out = 32'b00000000000000011011010011110100;
            12'b001100111011: out = 32'b00000000000000011011010110001011;
            12'b001100111100: out = 32'b00000000000000011011011000100010;
            12'b001100111101: out = 32'b00000000000000011011011010111010;
            12'b001100111110: out = 32'b00000000000000011011011101010001;
            12'b001100111111: out = 32'b00000000000000011011011111101001;
            12'b001101000000: out = 32'b00000000000000011011100010000001;
            12'b001101000001: out = 32'b00000000000000011011100100011000;
            12'b001101000010: out = 32'b00000000000000011011100110110000;
            12'b001101000011: out = 32'b00000000000000011011101001001000;
            12'b001101000100: out = 32'b00000000000000011011101011100000;
            12'b001101000101: out = 32'b00000000000000011011101101111000;
            12'b001101000110: out = 32'b00000000000000011011110000010000;
            12'b001101000111: out = 32'b00000000000000011011110010101000;
            12'b001101001000: out = 32'b00000000000000011011110101000000;
            12'b001101001001: out = 32'b00000000000000011011110111011000;
            12'b001101001010: out = 32'b00000000000000011011111001110001;
            12'b001101001011: out = 32'b00000000000000011011111100001001;
            12'b001101001100: out = 32'b00000000000000011011111110100001;
            12'b001101001101: out = 32'b00000000000000011100000000111010;
            12'b001101001110: out = 32'b00000000000000011100000011010011;
            12'b001101001111: out = 32'b00000000000000011100000101101011;
            12'b001101010000: out = 32'b00000000000000011100001000000100;
            12'b001101010001: out = 32'b00000000000000011100001010011101;
            12'b001101010010: out = 32'b00000000000000011100001100110101;
            12'b001101010011: out = 32'b00000000000000011100001111001110;
            12'b001101010100: out = 32'b00000000000000011100010001100111;
            12'b001101010101: out = 32'b00000000000000011100010100000000;
            12'b001101010110: out = 32'b00000000000000011100010110011001;
            12'b001101010111: out = 32'b00000000000000011100011000110011;
            12'b001101011000: out = 32'b00000000000000011100011011001100;
            12'b001101011001: out = 32'b00000000000000011100011101100101;
            12'b001101011010: out = 32'b00000000000000011100011111111110;
            12'b001101011011: out = 32'b00000000000000011100100010011000;
            12'b001101011100: out = 32'b00000000000000011100100100110001;
            12'b001101011101: out = 32'b00000000000000011100100111001011;
            12'b001101011110: out = 32'b00000000000000011100101001100100;
            12'b001101011111: out = 32'b00000000000000011100101011111110;
            12'b001101100000: out = 32'b00000000000000011100101110011000;
            12'b001101100001: out = 32'b00000000000000011100110000110010;
            12'b001101100010: out = 32'b00000000000000011100110011001100;
            12'b001101100011: out = 32'b00000000000000011100110101100110;
            12'b001101100100: out = 32'b00000000000000011100111000000000;
            12'b001101100101: out = 32'b00000000000000011100111010011010;
            12'b001101100110: out = 32'b00000000000000011100111100110100;
            12'b001101100111: out = 32'b00000000000000011100111111001110;
            12'b001101101000: out = 32'b00000000000000011101000001101000;
            12'b001101101001: out = 32'b00000000000000011101000100000011;
            12'b001101101010: out = 32'b00000000000000011101000110011101;
            12'b001101101011: out = 32'b00000000000000011101001000111000;
            12'b001101101100: out = 32'b00000000000000011101001011010010;
            12'b001101101101: out = 32'b00000000000000011101001101101101;
            12'b001101101110: out = 32'b00000000000000011101010000000111;
            12'b001101101111: out = 32'b00000000000000011101010010100010;
            12'b001101110000: out = 32'b00000000000000011101010100111101;
            12'b001101110001: out = 32'b00000000000000011101010111011000;
            12'b001101110010: out = 32'b00000000000000011101011001110011;
            12'b001101110011: out = 32'b00000000000000011101011100001110;
            12'b001101110100: out = 32'b00000000000000011101011110101001;
            12'b001101110101: out = 32'b00000000000000011101100001000100;
            12'b001101110110: out = 32'b00000000000000011101100011100000;
            12'b001101110111: out = 32'b00000000000000011101100101111011;
            12'b001101111000: out = 32'b00000000000000011101101000010110;
            12'b001101111001: out = 32'b00000000000000011101101010110010;
            12'b001101111010: out = 32'b00000000000000011101101101001101;
            12'b001101111011: out = 32'b00000000000000011101101111101001;
            12'b001101111100: out = 32'b00000000000000011101110010000101;
            12'b001101111101: out = 32'b00000000000000011101110100100000;
            12'b001101111110: out = 32'b00000000000000011101110110111100;
            12'b001101111111: out = 32'b00000000000000011101111001011000;
            12'b001110000000: out = 32'b00000000000000011101111011110100;
            12'b001110000001: out = 32'b00000000000000011101111110010000;
            12'b001110000010: out = 32'b00000000000000011110000000101100;
            12'b001110000011: out = 32'b00000000000000011110000011001000;
            12'b001110000100: out = 32'b00000000000000011110000101100101;
            12'b001110000101: out = 32'b00000000000000011110001000000001;
            12'b001110000110: out = 32'b00000000000000011110001010011101;
            12'b001110000111: out = 32'b00000000000000011110001100111010;
            12'b001110001000: out = 32'b00000000000000011110001111010110;
            12'b001110001001: out = 32'b00000000000000011110010001110011;
            12'b001110001010: out = 32'b00000000000000011110010100010000;
            12'b001110001011: out = 32'b00000000000000011110010110101100;
            12'b001110001100: out = 32'b00000000000000011110011001001001;
            12'b001110001101: out = 32'b00000000000000011110011011100110;
            12'b001110001110: out = 32'b00000000000000011110011110000011;
            12'b001110001111: out = 32'b00000000000000011110100000100000;
            12'b001110010000: out = 32'b00000000000000011110100010111101;
            12'b001110010001: out = 32'b00000000000000011110100101011011;
            12'b001110010010: out = 32'b00000000000000011110100111111000;
            12'b001110010011: out = 32'b00000000000000011110101010010101;
            12'b001110010100: out = 32'b00000000000000011110101100110011;
            12'b001110010101: out = 32'b00000000000000011110101111010000;
            12'b001110010110: out = 32'b00000000000000011110110001101110;
            12'b001110010111: out = 32'b00000000000000011110110100001011;
            12'b001110011000: out = 32'b00000000000000011110110110101001;
            12'b001110011001: out = 32'b00000000000000011110111001000111;
            12'b001110011010: out = 32'b00000000000000011110111011100101;
            12'b001110011011: out = 32'b00000000000000011110111110000011;
            12'b001110011100: out = 32'b00000000000000011111000000100001;
            12'b001110011101: out = 32'b00000000000000011111000010111111;
            12'b001110011110: out = 32'b00000000000000011111000101011101;
            12'b001110011111: out = 32'b00000000000000011111000111111011;
            12'b001110100000: out = 32'b00000000000000011111001010011001;
            12'b001110100001: out = 32'b00000000000000011111001100111000;
            12'b001110100010: out = 32'b00000000000000011111001111010110;
            12'b001110100011: out = 32'b00000000000000011111010001110101;
            12'b001110100100: out = 32'b00000000000000011111010100010011;
            12'b001110100101: out = 32'b00000000000000011111010110110010;
            12'b001110100110: out = 32'b00000000000000011111011001010001;
            12'b001110100111: out = 32'b00000000000000011111011011110000;
            12'b001110101000: out = 32'b00000000000000011111011110001111;
            12'b001110101001: out = 32'b00000000000000011111100000101110;
            12'b001110101010: out = 32'b00000000000000011111100011001101;
            12'b001110101011: out = 32'b00000000000000011111100101101100;
            12'b001110101100: out = 32'b00000000000000011111101000001011;
            12'b001110101101: out = 32'b00000000000000011111101010101010;
            12'b001110101110: out = 32'b00000000000000011111101101001010;
            12'b001110101111: out = 32'b00000000000000011111101111101001;
            12'b001110110000: out = 32'b00000000000000011111110010001001;
            12'b001110110001: out = 32'b00000000000000011111110100101000;
            12'b001110110010: out = 32'b00000000000000011111110111001000;
            12'b001110110011: out = 32'b00000000000000011111111001101000;
            12'b001110110100: out = 32'b00000000000000011111111100001000;
            12'b001110110101: out = 32'b00000000000000011111111110100111;
            12'b001110110110: out = 32'b00000000000000100000000001000111;
            12'b001110110111: out = 32'b00000000000000100000000011101000;
            12'b001110111000: out = 32'b00000000000000100000000110001000;
            12'b001110111001: out = 32'b00000000000000100000001000101000;
            12'b001110111010: out = 32'b00000000000000100000001011001000;
            12'b001110111011: out = 32'b00000000000000100000001101101001;
            12'b001110111100: out = 32'b00000000000000100000010000001001;
            12'b001110111101: out = 32'b00000000000000100000010010101010;
            12'b001110111110: out = 32'b00000000000000100000010101001010;
            12'b001110111111: out = 32'b00000000000000100000010111101011;
            12'b001111000000: out = 32'b00000000000000100000011010001100;
            12'b001111000001: out = 32'b00000000000000100000011100101101;
            12'b001111000010: out = 32'b00000000000000100000011111001110;
            12'b001111000011: out = 32'b00000000000000100000100001101111;
            12'b001111000100: out = 32'b00000000000000100000100100010000;
            12'b001111000101: out = 32'b00000000000000100000100110110001;
            12'b001111000110: out = 32'b00000000000000100000101001010010;
            12'b001111000111: out = 32'b00000000000000100000101011110011;
            12'b001111001000: out = 32'b00000000000000100000101110010101;
            12'b001111001001: out = 32'b00000000000000100000110000110110;
            12'b001111001010: out = 32'b00000000000000100000110011011000;
            12'b001111001011: out = 32'b00000000000000100000110101111010;
            12'b001111001100: out = 32'b00000000000000100000111000011011;
            12'b001111001101: out = 32'b00000000000000100000111010111101;
            12'b001111001110: out = 32'b00000000000000100000111101011111;
            12'b001111001111: out = 32'b00000000000000100001000000000001;
            12'b001111010000: out = 32'b00000000000000100001000010100011;
            12'b001111010001: out = 32'b00000000000000100001000101000101;
            12'b001111010010: out = 32'b00000000000000100001000111101000;
            12'b001111010011: out = 32'b00000000000000100001001010001010;
            12'b001111010100: out = 32'b00000000000000100001001100101100;
            12'b001111010101: out = 32'b00000000000000100001001111001111;
            12'b001111010110: out = 32'b00000000000000100001010001110001;
            12'b001111010111: out = 32'b00000000000000100001010100010100;
            12'b001111011000: out = 32'b00000000000000100001010110110111;
            12'b001111011001: out = 32'b00000000000000100001011001011010;
            12'b001111011010: out = 32'b00000000000000100001011011111100;
            12'b001111011011: out = 32'b00000000000000100001011110011111;
            12'b001111011100: out = 32'b00000000000000100001100001000010;
            12'b001111011101: out = 32'b00000000000000100001100011100110;
            12'b001111011110: out = 32'b00000000000000100001100110001001;
            12'b001111011111: out = 32'b00000000000000100001101000101100;
            12'b001111100000: out = 32'b00000000000000100001101011010000;
            12'b001111100001: out = 32'b00000000000000100001101101110011;
            12'b001111100010: out = 32'b00000000000000100001110000010111;
            12'b001111100011: out = 32'b00000000000000100001110010111010;
            12'b001111100100: out = 32'b00000000000000100001110101011110;
            12'b001111100101: out = 32'b00000000000000100001111000000010;
            12'b001111100110: out = 32'b00000000000000100001111010100110;
            12'b001111100111: out = 32'b00000000000000100001111101001010;
            12'b001111101000: out = 32'b00000000000000100001111111101110;
            12'b001111101001: out = 32'b00000000000000100010000010010010;
            12'b001111101010: out = 32'b00000000000000100010000100110110;
            12'b001111101011: out = 32'b00000000000000100010000111011011;
            12'b001111101100: out = 32'b00000000000000100010001001111111;
            12'b001111101101: out = 32'b00000000000000100010001100100011;
            12'b001111101110: out = 32'b00000000000000100010001111001000;
            12'b001111101111: out = 32'b00000000000000100010010001101101;
            12'b001111110000: out = 32'b00000000000000100010010100010001;
            12'b001111110001: out = 32'b00000000000000100010010110110110;
            12'b001111110010: out = 32'b00000000000000100010011001011011;
            12'b001111110011: out = 32'b00000000000000100010011100000000;
            12'b001111110100: out = 32'b00000000000000100010011110100101;
            12'b001111110101: out = 32'b00000000000000100010100001001011;
            12'b001111110110: out = 32'b00000000000000100010100011110000;
            12'b001111110111: out = 32'b00000000000000100010100110010101;
            12'b001111111000: out = 32'b00000000000000100010101000111011;
            12'b001111111001: out = 32'b00000000000000100010101011100000;
            12'b001111111010: out = 32'b00000000000000100010101110000110;
            12'b001111111011: out = 32'b00000000000000100010110000101100;
            12'b001111111100: out = 32'b00000000000000100010110011010001;
            12'b001111111101: out = 32'b00000000000000100010110101110111;
            12'b001111111110: out = 32'b00000000000000100010111000011101;
            12'b001111111111: out = 32'b00000000000000100010111011000011;
            12'b010000000000: out = 32'b00000000000000100010111101101001;
            12'b010000000001: out = 32'b00000000000000100011000000010000;
            12'b010000000010: out = 32'b00000000000000100011000010110110;
            12'b010000000011: out = 32'b00000000000000100011000101011100;
            12'b010000000100: out = 32'b00000000000000100011001000000011;
            12'b010000000101: out = 32'b00000000000000100011001010101010;
            12'b010000000110: out = 32'b00000000000000100011001101010000;
            12'b010000000111: out = 32'b00000000000000100011001111110111;
            12'b010000001000: out = 32'b00000000000000100011010010011110;
            12'b010000001001: out = 32'b00000000000000100011010101000101;
            12'b010000001010: out = 32'b00000000000000100011010111101100;
            12'b010000001011: out = 32'b00000000000000100011011010010011;
            12'b010000001100: out = 32'b00000000000000100011011100111010;
            12'b010000001101: out = 32'b00000000000000100011011111100010;
            12'b010000001110: out = 32'b00000000000000100011100010001001;
            12'b010000001111: out = 32'b00000000000000100011100100110000;
            12'b010000010000: out = 32'b00000000000000100011100111011000;
            12'b010000010001: out = 32'b00000000000000100011101010000000;
            12'b010000010010: out = 32'b00000000000000100011101100101000;
            12'b010000010011: out = 32'b00000000000000100011101111001111;
            12'b010000010100: out = 32'b00000000000000100011110001110111;
            12'b010000010101: out = 32'b00000000000000100011110100011111;
            12'b010000010110: out = 32'b00000000000000100011110111001000;
            12'b010000010111: out = 32'b00000000000000100011111001110000;
            12'b010000011000: out = 32'b00000000000000100011111100011000;
            12'b010000011001: out = 32'b00000000000000100011111111000001;
            12'b010000011010: out = 32'b00000000000000100100000001101001;
            12'b010000011011: out = 32'b00000000000000100100000100010010;
            12'b010000011100: out = 32'b00000000000000100100000110111010;
            12'b010000011101: out = 32'b00000000000000100100001001100011;
            12'b010000011110: out = 32'b00000000000000100100001100001100;
            12'b010000011111: out = 32'b00000000000000100100001110110101;
            12'b010000100000: out = 32'b00000000000000100100010001011110;
            12'b010000100001: out = 32'b00000000000000100100010100000111;
            12'b010000100010: out = 32'b00000000000000100100010110110001;
            12'b010000100011: out = 32'b00000000000000100100011001011010;
            12'b010000100100: out = 32'b00000000000000100100011100000011;
            12'b010000100101: out = 32'b00000000000000100100011110101101;
            12'b010000100110: out = 32'b00000000000000100100100001010110;
            12'b010000100111: out = 32'b00000000000000100100100100000000;
            12'b010000101000: out = 32'b00000000000000100100100110101010;
            12'b010000101001: out = 32'b00000000000000100100101001010100;
            12'b010000101010: out = 32'b00000000000000100100101011111110;
            12'b010000101011: out = 32'b00000000000000100100101110101000;
            12'b010000101100: out = 32'b00000000000000100100110001010010;
            12'b010000101101: out = 32'b00000000000000100100110011111101;
            12'b010000101110: out = 32'b00000000000000100100110110100111;
            12'b010000101111: out = 32'b00000000000000100100111001010001;
            12'b010000110000: out = 32'b00000000000000100100111011111100;
            12'b010000110001: out = 32'b00000000000000100100111110100111;
            12'b010000110010: out = 32'b00000000000000100101000001010010;
            12'b010000110011: out = 32'b00000000000000100101000011111100;
            12'b010000110100: out = 32'b00000000000000100101000110100111;
            12'b010000110101: out = 32'b00000000000000100101001001010010;
            12'b010000110110: out = 32'b00000000000000100101001011111110;
            12'b010000110111: out = 32'b00000000000000100101001110101001;
            12'b010000111000: out = 32'b00000000000000100101010001010100;
            12'b010000111001: out = 32'b00000000000000100101010100000000;
            12'b010000111010: out = 32'b00000000000000100101010110101011;
            12'b010000111011: out = 32'b00000000000000100101011001010111;
            12'b010000111100: out = 32'b00000000000000100101011100000011;
            12'b010000111101: out = 32'b00000000000000100101011110101110;
            12'b010000111110: out = 32'b00000000000000100101100001011010;
            12'b010000111111: out = 32'b00000000000000100101100100000110;
            12'b010001000000: out = 32'b00000000000000100101100110110011;
            12'b010001000001: out = 32'b00000000000000100101101001011111;
            12'b010001000010: out = 32'b00000000000000100101101100001011;
            12'b010001000011: out = 32'b00000000000000100101101110111000;
            12'b010001000100: out = 32'b00000000000000100101110001100100;
            12'b010001000101: out = 32'b00000000000000100101110100010001;
            12'b010001000110: out = 32'b00000000000000100101110110111110;
            12'b010001000111: out = 32'b00000000000000100101111001101010;
            12'b010001001000: out = 32'b00000000000000100101111100010111;
            12'b010001001001: out = 32'b00000000000000100101111111000100;
            12'b010001001010: out = 32'b00000000000000100110000001110010;
            12'b010001001011: out = 32'b00000000000000100110000100011111;
            12'b010001001100: out = 32'b00000000000000100110000111001100;
            12'b010001001101: out = 32'b00000000000000100110001001111010;
            12'b010001001110: out = 32'b00000000000000100110001100100111;
            12'b010001001111: out = 32'b00000000000000100110001111010101;
            12'b010001010000: out = 32'b00000000000000100110010010000011;
            12'b010001010001: out = 32'b00000000000000100110010100110000;
            12'b010001010010: out = 32'b00000000000000100110010111011110;
            12'b010001010011: out = 32'b00000000000000100110011010001100;
            12'b010001010100: out = 32'b00000000000000100110011100111011;
            12'b010001010101: out = 32'b00000000000000100110011111101001;
            12'b010001010110: out = 32'b00000000000000100110100010010111;
            12'b010001010111: out = 32'b00000000000000100110100101000110;
            12'b010001011000: out = 32'b00000000000000100110100111110100;
            12'b010001011001: out = 32'b00000000000000100110101010100011;
            12'b010001011010: out = 32'b00000000000000100110101101010010;
            12'b010001011011: out = 32'b00000000000000100110110000000000;
            12'b010001011100: out = 32'b00000000000000100110110010101111;
            12'b010001011101: out = 32'b00000000000000100110110101011111;
            12'b010001011110: out = 32'b00000000000000100110111000001110;
            12'b010001011111: out = 32'b00000000000000100110111010111101;
            12'b010001100000: out = 32'b00000000000000100110111101101100;
            12'b010001100001: out = 32'b00000000000000100111000000011100;
            12'b010001100010: out = 32'b00000000000000100111000011001011;
            12'b010001100011: out = 32'b00000000000000100111000101111011;
            12'b010001100100: out = 32'b00000000000000100111001000101011;
            12'b010001100101: out = 32'b00000000000000100111001011011011;
            12'b010001100110: out = 32'b00000000000000100111001110001011;
            12'b010001100111: out = 32'b00000000000000100111010000111011;
            12'b010001101000: out = 32'b00000000000000100111010011101011;
            12'b010001101001: out = 32'b00000000000000100111010110011100;
            12'b010001101010: out = 32'b00000000000000100111011001001100;
            12'b010001101011: out = 32'b00000000000000100111011011111101;
            12'b010001101100: out = 32'b00000000000000100111011110101101;
            12'b010001101101: out = 32'b00000000000000100111100001011110;
            12'b010001101110: out = 32'b00000000000000100111100100001111;
            12'b010001101111: out = 32'b00000000000000100111100111000000;
            12'b010001110000: out = 32'b00000000000000100111101001110001;
            12'b010001110001: out = 32'b00000000000000100111101100100010;
            12'b010001110010: out = 32'b00000000000000100111101111010011;
            12'b010001110011: out = 32'b00000000000000100111110010000101;
            12'b010001110100: out = 32'b00000000000000100111110100110110;
            12'b010001110101: out = 32'b00000000000000100111110111101000;
            12'b010001110110: out = 32'b00000000000000100111111010011010;
            12'b010001110111: out = 32'b00000000000000100111111101001100;
            12'b010001111000: out = 32'b00000000000000100111111111111101;
            12'b010001111001: out = 32'b00000000000000101000000010110000;
            12'b010001111010: out = 32'b00000000000000101000000101100010;
            12'b010001111011: out = 32'b00000000000000101000001000010100;
            12'b010001111100: out = 32'b00000000000000101000001011000110;
            12'b010001111101: out = 32'b00000000000000101000001101111001;
            12'b010001111110: out = 32'b00000000000000101000010000101011;
            12'b010001111111: out = 32'b00000000000000101000010011011110;
            12'b010010000000: out = 32'b00000000000000101000010110010001;
            12'b010010000001: out = 32'b00000000000000101000011001000100;
            12'b010010000010: out = 32'b00000000000000101000011011110111;
            12'b010010000011: out = 32'b00000000000000101000011110101010;
            12'b010010000100: out = 32'b00000000000000101000100001011101;
            12'b010010000101: out = 32'b00000000000000101000100100010001;
            12'b010010000110: out = 32'b00000000000000101000100111000100;
            12'b010010000111: out = 32'b00000000000000101000101001111000;
            12'b010010001000: out = 32'b00000000000000101000101100101011;
            12'b010010001001: out = 32'b00000000000000101000101111011111;
            12'b010010001010: out = 32'b00000000000000101000110010010011;
            12'b010010001011: out = 32'b00000000000000101000110101000111;
            12'b010010001100: out = 32'b00000000000000101000110111111011;
            12'b010010001101: out = 32'b00000000000000101000111010110000;
            12'b010010001110: out = 32'b00000000000000101000111101100100;
            12'b010010001111: out = 32'b00000000000000101001000000011001;
            12'b010010010000: out = 32'b00000000000000101001000011001101;
            12'b010010010001: out = 32'b00000000000000101001000110000010;
            12'b010010010010: out = 32'b00000000000000101001001000110111;
            12'b010010010011: out = 32'b00000000000000101001001011101100;
            12'b010010010100: out = 32'b00000000000000101001001110100001;
            12'b010010010101: out = 32'b00000000000000101001010001010110;
            12'b010010010110: out = 32'b00000000000000101001010100001011;
            12'b010010010111: out = 32'b00000000000000101001010111000001;
            12'b010010011000: out = 32'b00000000000000101001011001110110;
            12'b010010011001: out = 32'b00000000000000101001011100101100;
            12'b010010011010: out = 32'b00000000000000101001011111100001;
            12'b010010011011: out = 32'b00000000000000101001100010010111;
            12'b010010011100: out = 32'b00000000000000101001100101001101;
            12'b010010011101: out = 32'b00000000000000101001101000000011;
            12'b010010011110: out = 32'b00000000000000101001101010111010;
            12'b010010011111: out = 32'b00000000000000101001101101110000;
            12'b010010100000: out = 32'b00000000000000101001110000100110;
            12'b010010100001: out = 32'b00000000000000101001110011011101;
            12'b010010100010: out = 32'b00000000000000101001110110010100;
            12'b010010100011: out = 32'b00000000000000101001111001001010;
            12'b010010100100: out = 32'b00000000000000101001111100000001;
            12'b010010100101: out = 32'b00000000000000101001111110111000;
            12'b010010100110: out = 32'b00000000000000101010000001101111;
            12'b010010100111: out = 32'b00000000000000101010000100100111;
            12'b010010101000: out = 32'b00000000000000101010000111011110;
            12'b010010101001: out = 32'b00000000000000101010001010010110;
            12'b010010101010: out = 32'b00000000000000101010001101001101;
            12'b010010101011: out = 32'b00000000000000101010010000000101;
            12'b010010101100: out = 32'b00000000000000101010010010111101;
            12'b010010101101: out = 32'b00000000000000101010010101110101;
            12'b010010101110: out = 32'b00000000000000101010011000101101;
            12'b010010101111: out = 32'b00000000000000101010011011100101;
            12'b010010110000: out = 32'b00000000000000101010011110011101;
            12'b010010110001: out = 32'b00000000000000101010100001010110;
            12'b010010110010: out = 32'b00000000000000101010100100001110;
            12'b010010110011: out = 32'b00000000000000101010100111000111;
            12'b010010110100: out = 32'b00000000000000101010101010000000;
            12'b010010110101: out = 32'b00000000000000101010101100111001;
            12'b010010110110: out = 32'b00000000000000101010101111110010;
            12'b010010110111: out = 32'b00000000000000101010110010101011;
            12'b010010111000: out = 32'b00000000000000101010110101100100;
            12'b010010111001: out = 32'b00000000000000101010111000011110;
            12'b010010111010: out = 32'b00000000000000101010111011010111;
            12'b010010111011: out = 32'b00000000000000101010111110010001;
            12'b010010111100: out = 32'b00000000000000101011000001001011;
            12'b010010111101: out = 32'b00000000000000101011000100000100;
            12'b010010111110: out = 32'b00000000000000101011000110111110;
            12'b010010111111: out = 32'b00000000000000101011001001111001;
            12'b010011000000: out = 32'b00000000000000101011001100110011;
            12'b010011000001: out = 32'b00000000000000101011001111101101;
            12'b010011000010: out = 32'b00000000000000101011010010101000;
            12'b010011000011: out = 32'b00000000000000101011010101100010;
            12'b010011000100: out = 32'b00000000000000101011011000011101;
            12'b010011000101: out = 32'b00000000000000101011011011011000;
            12'b010011000110: out = 32'b00000000000000101011011110010011;
            12'b010011000111: out = 32'b00000000000000101011100001001110;
            12'b010011001000: out = 32'b00000000000000101011100100001001;
            12'b010011001001: out = 32'b00000000000000101011100111000101;
            12'b010011001010: out = 32'b00000000000000101011101010000000;
            12'b010011001011: out = 32'b00000000000000101011101100111100;
            12'b010011001100: out = 32'b00000000000000101011101111111000;
            12'b010011001101: out = 32'b00000000000000101011110010110011;
            12'b010011001110: out = 32'b00000000000000101011110101101111;
            12'b010011001111: out = 32'b00000000000000101011111000101100;
            12'b010011010000: out = 32'b00000000000000101011111011101000;
            12'b010011010001: out = 32'b00000000000000101011111110100100;
            12'b010011010010: out = 32'b00000000000000101100000001100001;
            12'b010011010011: out = 32'b00000000000000101100000100011101;
            12'b010011010100: out = 32'b00000000000000101100000111011010;
            12'b010011010101: out = 32'b00000000000000101100001010010111;
            12'b010011010110: out = 32'b00000000000000101100001101010100;
            12'b010011010111: out = 32'b00000000000000101100010000010001;
            12'b010011011000: out = 32'b00000000000000101100010011001110;
            12'b010011011001: out = 32'b00000000000000101100010110001100;
            12'b010011011010: out = 32'b00000000000000101100011001001001;
            12'b010011011011: out = 32'b00000000000000101100011100000111;
            12'b010011011100: out = 32'b00000000000000101100011111000101;
            12'b010011011101: out = 32'b00000000000000101100100010000011;
            12'b010011011110: out = 32'b00000000000000101100100101000001;
            12'b010011011111: out = 32'b00000000000000101100100111111111;
            12'b010011100000: out = 32'b00000000000000101100101010111101;
            12'b010011100001: out = 32'b00000000000000101100101101111100;
            12'b010011100010: out = 32'b00000000000000101100110000111010;
            12'b010011100011: out = 32'b00000000000000101100110011111001;
            12'b010011100100: out = 32'b00000000000000101100110110111000;
            12'b010011100101: out = 32'b00000000000000101100111001110111;
            12'b010011100110: out = 32'b00000000000000101100111100110110;
            12'b010011100111: out = 32'b00000000000000101100111111110101;
            12'b010011101000: out = 32'b00000000000000101101000010110100;
            12'b010011101001: out = 32'b00000000000000101101000101110100;
            12'b010011101010: out = 32'b00000000000000101101001000110011;
            12'b010011101011: out = 32'b00000000000000101101001011110011;
            12'b010011101100: out = 32'b00000000000000101101001110110011;
            12'b010011101101: out = 32'b00000000000000101101010001110011;
            12'b010011101110: out = 32'b00000000000000101101010100110011;
            12'b010011101111: out = 32'b00000000000000101101010111110011;
            12'b010011110000: out = 32'b00000000000000101101011010110100;
            12'b010011110001: out = 32'b00000000000000101101011101110100;
            12'b010011110010: out = 32'b00000000000000101101100000110101;
            12'b010011110011: out = 32'b00000000000000101101100011110110;
            12'b010011110100: out = 32'b00000000000000101101100110110111;
            12'b010011110101: out = 32'b00000000000000101101101001111000;
            12'b010011110110: out = 32'b00000000000000101101101100111001;
            12'b010011110111: out = 32'b00000000000000101101101111111010;
            12'b010011111000: out = 32'b00000000000000101101110010111100;
            12'b010011111001: out = 32'b00000000000000101101110101111101;
            12'b010011111010: out = 32'b00000000000000101101111000111111;
            12'b010011111011: out = 32'b00000000000000101101111100000001;
            12'b010011111100: out = 32'b00000000000000101101111111000011;
            12'b010011111101: out = 32'b00000000000000101110000010000101;
            12'b010011111110: out = 32'b00000000000000101110000101000111;
            12'b010011111111: out = 32'b00000000000000101110001000001010;
            12'b010100000000: out = 32'b00000000000000101110001011001100;
            12'b010100000001: out = 32'b00000000000000101110001110001111;
            12'b010100000010: out = 32'b00000000000000101110010001010010;
            12'b010100000011: out = 32'b00000000000000101110010100010101;
            12'b010100000100: out = 32'b00000000000000101110010111011000;
            12'b010100000101: out = 32'b00000000000000101110011010011011;
            12'b010100000110: out = 32'b00000000000000101110011101011111;
            12'b010100000111: out = 32'b00000000000000101110100000100010;
            12'b010100001000: out = 32'b00000000000000101110100011100110;
            12'b010100001001: out = 32'b00000000000000101110100110101010;
            12'b010100001010: out = 32'b00000000000000101110101001101110;
            12'b010100001011: out = 32'b00000000000000101110101100110010;
            12'b010100001100: out = 32'b00000000000000101110101111110110;
            12'b010100001101: out = 32'b00000000000000101110110010111010;
            12'b010100001110: out = 32'b00000000000000101110110101111111;
            12'b010100001111: out = 32'b00000000000000101110111001000011;
            12'b010100010000: out = 32'b00000000000000101110111100001000;
            12'b010100010001: out = 32'b00000000000000101110111111001101;
            12'b010100010010: out = 32'b00000000000000101111000010010010;
            12'b010100010011: out = 32'b00000000000000101111000101010111;
            12'b010100010100: out = 32'b00000000000000101111001000011101;
            12'b010100010101: out = 32'b00000000000000101111001011100010;
            12'b010100010110: out = 32'b00000000000000101111001110101000;
            12'b010100010111: out = 32'b00000000000000101111010001101110;
            12'b010100011000: out = 32'b00000000000000101111010100110011;
            12'b010100011001: out = 32'b00000000000000101111010111111010;
            12'b010100011010: out = 32'b00000000000000101111011011000000;
            12'b010100011011: out = 32'b00000000000000101111011110000110;
            12'b010100011100: out = 32'b00000000000000101111100001001101;
            12'b010100011101: out = 32'b00000000000000101111100100010011;
            12'b010100011110: out = 32'b00000000000000101111100111011010;
            12'b010100011111: out = 32'b00000000000000101111101010100001;
            12'b010100100000: out = 32'b00000000000000101111101101101000;
            12'b010100100001: out = 32'b00000000000000101111110000101111;
            12'b010100100010: out = 32'b00000000000000101111110011110111;
            12'b010100100011: out = 32'b00000000000000101111110110111110;
            12'b010100100100: out = 32'b00000000000000101111111010000110;
            12'b010100100101: out = 32'b00000000000000101111111101001110;
            12'b010100100110: out = 32'b00000000000000110000000000010101;
            12'b010100100111: out = 32'b00000000000000110000000011011110;
            12'b010100101000: out = 32'b00000000000000110000000110100110;
            12'b010100101001: out = 32'b00000000000000110000001001101110;
            12'b010100101010: out = 32'b00000000000000110000001100110111;
            12'b010100101011: out = 32'b00000000000000110000001111111111;
            12'b010100101100: out = 32'b00000000000000110000010011001000;
            12'b010100101101: out = 32'b00000000000000110000010110010001;
            12'b010100101110: out = 32'b00000000000000110000011001011010;
            12'b010100101111: out = 32'b00000000000000110000011100100100;
            12'b010100110000: out = 32'b00000000000000110000011111101101;
            12'b010100110001: out = 32'b00000000000000110000100010110111;
            12'b010100110010: out = 32'b00000000000000110000100110000000;
            12'b010100110011: out = 32'b00000000000000110000101001001010;
            12'b010100110100: out = 32'b00000000000000110000101100010100;
            12'b010100110101: out = 32'b00000000000000110000101111011110;
            12'b010100110110: out = 32'b00000000000000110000110010101001;
            12'b010100110111: out = 32'b00000000000000110000110101110011;
            12'b010100111000: out = 32'b00000000000000110000111000111110;
            12'b010100111001: out = 32'b00000000000000110000111100001000;
            12'b010100111010: out = 32'b00000000000000110000111111010011;
            12'b010100111011: out = 32'b00000000000000110001000010011110;
            12'b010100111100: out = 32'b00000000000000110001000101101010;
            12'b010100111101: out = 32'b00000000000000110001001000110101;
            12'b010100111110: out = 32'b00000000000000110001001100000001;
            12'b010100111111: out = 32'b00000000000000110001001111001100;
            12'b010101000000: out = 32'b00000000000000110001010010011000;
            12'b010101000001: out = 32'b00000000000000110001010101100100;
            12'b010101000010: out = 32'b00000000000000110001011000110000;
            12'b010101000011: out = 32'b00000000000000110001011011111101;
            12'b010101000100: out = 32'b00000000000000110001011111001001;
            12'b010101000101: out = 32'b00000000000000110001100010010110;
            12'b010101000110: out = 32'b00000000000000110001100101100010;
            12'b010101000111: out = 32'b00000000000000110001101000101111;
            12'b010101001000: out = 32'b00000000000000110001101011111100;
            12'b010101001001: out = 32'b00000000000000110001101111001010;
            12'b010101001010: out = 32'b00000000000000110001110010010111;
            12'b010101001011: out = 32'b00000000000000110001110101100101;
            12'b010101001100: out = 32'b00000000000000110001111000110010;
            12'b010101001101: out = 32'b00000000000000110001111100000000;
            12'b010101001110: out = 32'b00000000000000110001111111001110;
            12'b010101001111: out = 32'b00000000000000110010000010011100;
            12'b010101010000: out = 32'b00000000000000110010000101101011;
            12'b010101010001: out = 32'b00000000000000110010001000111001;
            12'b010101010010: out = 32'b00000000000000110010001100001000;
            12'b010101010011: out = 32'b00000000000000110010001111010110;
            12'b010101010100: out = 32'b00000000000000110010010010100101;
            12'b010101010101: out = 32'b00000000000000110010010101110101;
            12'b010101010110: out = 32'b00000000000000110010011001000100;
            12'b010101010111: out = 32'b00000000000000110010011100010011;
            12'b010101011000: out = 32'b00000000000000110010011111100011;
            12'b010101011001: out = 32'b00000000000000110010100010110011;
            12'b010101011010: out = 32'b00000000000000110010100110000011;
            12'b010101011011: out = 32'b00000000000000110010101001010011;
            12'b010101011100: out = 32'b00000000000000110010101100100011;
            12'b010101011101: out = 32'b00000000000000110010101111110011;
            12'b010101011110: out = 32'b00000000000000110010110011000100;
            12'b010101011111: out = 32'b00000000000000110010110110010101;
            12'b010101100000: out = 32'b00000000000000110010111001100101;
            12'b010101100001: out = 32'b00000000000000110010111100110110;
            12'b010101100010: out = 32'b00000000000000110011000000001000;
            12'b010101100011: out = 32'b00000000000000110011000011011001;
            12'b010101100100: out = 32'b00000000000000110011000110101011;
            12'b010101100101: out = 32'b00000000000000110011001001111100;
            12'b010101100110: out = 32'b00000000000000110011001101001110;
            12'b010101100111: out = 32'b00000000000000110011010000100000;
            12'b010101101000: out = 32'b00000000000000110011010011110010;
            12'b010101101001: out = 32'b00000000000000110011010111000101;
            12'b010101101010: out = 32'b00000000000000110011011010010111;
            12'b010101101011: out = 32'b00000000000000110011011101101010;
            12'b010101101100: out = 32'b00000000000000110011100000111101;
            12'b010101101101: out = 32'b00000000000000110011100100010000;
            12'b010101101110: out = 32'b00000000000000110011100111100011;
            12'b010101101111: out = 32'b00000000000000110011101010110110;
            12'b010101110000: out = 32'b00000000000000110011101110001010;
            12'b010101110001: out = 32'b00000000000000110011110001011101;
            12'b010101110010: out = 32'b00000000000000110011110100110001;
            12'b010101110011: out = 32'b00000000000000110011111000000101;
            12'b010101110100: out = 32'b00000000000000110011111011011001;
            12'b010101110101: out = 32'b00000000000000110011111110101110;
            12'b010101110110: out = 32'b00000000000000110100000010000010;
            12'b010101110111: out = 32'b00000000000000110100000101010111;
            12'b010101111000: out = 32'b00000000000000110100001000101100;
            12'b010101111001: out = 32'b00000000000000110100001100000001;
            12'b010101111010: out = 32'b00000000000000110100001111010110;
            12'b010101111011: out = 32'b00000000000000110100010010101100;
            12'b010101111100: out = 32'b00000000000000110100010110000001;
            12'b010101111101: out = 32'b00000000000000110100011001010111;
            12'b010101111110: out = 32'b00000000000000110100011100101101;
            12'b010101111111: out = 32'b00000000000000110100100000000011;
            12'b010110000000: out = 32'b00000000000000110100100011011001;
            12'b010110000001: out = 32'b00000000000000110100100110101111;
            12'b010110000010: out = 32'b00000000000000110100101010000110;
            12'b010110000011: out = 32'b00000000000000110100101101011101;
            12'b010110000100: out = 32'b00000000000000110100110000110100;
            12'b010110000101: out = 32'b00000000000000110100110100001011;
            12'b010110000110: out = 32'b00000000000000110100110111100010;
            12'b010110000111: out = 32'b00000000000000110100111010111001;
            12'b010110001000: out = 32'b00000000000000110100111110010001;
            12'b010110001001: out = 32'b00000000000000110101000001101001;
            12'b010110001010: out = 32'b00000000000000110101000101000001;
            12'b010110001011: out = 32'b00000000000000110101001000011001;
            12'b010110001100: out = 32'b00000000000000110101001011110001;
            12'b010110001101: out = 32'b00000000000000110101001111001010;
            12'b010110001110: out = 32'b00000000000000110101010010100010;
            12'b010110001111: out = 32'b00000000000000110101010101111011;
            12'b010110010000: out = 32'b00000000000000110101011001010100;
            12'b010110010001: out = 32'b00000000000000110101011100101101;
            12'b010110010010: out = 32'b00000000000000110101100000000111;
            12'b010110010011: out = 32'b00000000000000110101100011100000;
            12'b010110010100: out = 32'b00000000000000110101100110111010;
            12'b010110010101: out = 32'b00000000000000110101101010010100;
            12'b010110010110: out = 32'b00000000000000110101101101101110;
            12'b010110010111: out = 32'b00000000000000110101110001001000;
            12'b010110011000: out = 32'b00000000000000110101110100100010;
            12'b010110011001: out = 32'b00000000000000110101110111111101;
            12'b010110011010: out = 32'b00000000000000110101111011011000;
            12'b010110011011: out = 32'b00000000000000110101111110110011;
            12'b010110011100: out = 32'b00000000000000110110000010001110;
            12'b010110011101: out = 32'b00000000000000110110000101101001;
            12'b010110011110: out = 32'b00000000000000110110001001000101;
            12'b010110011111: out = 32'b00000000000000110110001100100001;
            12'b010110100000: out = 32'b00000000000000110110001111111100;
            12'b010110100001: out = 32'b00000000000000110110010011011000;
            12'b010110100010: out = 32'b00000000000000110110010110110101;
            12'b010110100011: out = 32'b00000000000000110110011010010001;
            12'b010110100100: out = 32'b00000000000000110110011101101110;
            12'b010110100101: out = 32'b00000000000000110110100001001011;
            12'b010110100110: out = 32'b00000000000000110110100100101000;
            12'b010110100111: out = 32'b00000000000000110110101000000101;
            12'b010110101000: out = 32'b00000000000000110110101011100010;
            12'b010110101001: out = 32'b00000000000000110110101111000000;
            12'b010110101010: out = 32'b00000000000000110110110010011101;
            12'b010110101011: out = 32'b00000000000000110110110101111011;
            12'b010110101100: out = 32'b00000000000000110110111001011001;
            12'b010110101101: out = 32'b00000000000000110110111100111000;
            12'b010110101110: out = 32'b00000000000000110111000000010110;
            12'b010110101111: out = 32'b00000000000000110111000011110101;
            12'b010110110000: out = 32'b00000000000000110111000111010011;
            12'b010110110001: out = 32'b00000000000000110111001010110010;
            12'b010110110010: out = 32'b00000000000000110111001110010010;
            12'b010110110011: out = 32'b00000000000000110111010001110001;
            12'b010110110100: out = 32'b00000000000000110111010101010001;
            12'b010110110101: out = 32'b00000000000000110111011000110000;
            12'b010110110110: out = 32'b00000000000000110111011100010000;
            12'b010110110111: out = 32'b00000000000000110111011111110001;
            12'b010110111000: out = 32'b00000000000000110111100011010001;
            12'b010110111001: out = 32'b00000000000000110111100110110001;
            12'b010110111010: out = 32'b00000000000000110111101010010010;
            12'b010110111011: out = 32'b00000000000000110111101101110011;
            12'b010110111100: out = 32'b00000000000000110111110001010100;
            12'b010110111101: out = 32'b00000000000000110111110100110101;
            12'b010110111110: out = 32'b00000000000000110111111000010111;
            12'b010110111111: out = 32'b00000000000000110111111011111001;
            12'b010111000000: out = 32'b00000000000000110111111111011010;
            12'b010111000001: out = 32'b00000000000000111000000010111101;
            12'b010111000010: out = 32'b00000000000000111000000110011111;
            12'b010111000011: out = 32'b00000000000000111000001010000001;
            12'b010111000100: out = 32'b00000000000000111000001101100100;
            12'b010111000101: out = 32'b00000000000000111000010001000111;
            12'b010111000110: out = 32'b00000000000000111000010100101010;
            12'b010111000111: out = 32'b00000000000000111000011000001101;
            12'b010111001000: out = 32'b00000000000000111000011011110000;
            12'b010111001001: out = 32'b00000000000000111000011111010100;
            12'b010111001010: out = 32'b00000000000000111000100010111000;
            12'b010111001011: out = 32'b00000000000000111000100110011100;
            12'b010111001100: out = 32'b00000000000000111000101010000000;
            12'b010111001101: out = 32'b00000000000000111000101101100101;
            12'b010111001110: out = 32'b00000000000000111000110001001001;
            12'b010111001111: out = 32'b00000000000000111000110100101110;
            12'b010111010000: out = 32'b00000000000000111000111000010011;
            12'b010111010001: out = 32'b00000000000000111000111011111000;
            12'b010111010010: out = 32'b00000000000000111000111111011110;
            12'b010111010011: out = 32'b00000000000000111001000011000011;
            12'b010111010100: out = 32'b00000000000000111001000110101001;
            12'b010111010101: out = 32'b00000000000000111001001010001111;
            12'b010111010110: out = 32'b00000000000000111001001101110101;
            12'b010111010111: out = 32'b00000000000000111001010001011100;
            12'b010111011000: out = 32'b00000000000000111001010101000010;
            12'b010111011001: out = 32'b00000000000000111001011000101001;
            12'b010111011010: out = 32'b00000000000000111001011100010000;
            12'b010111011011: out = 32'b00000000000000111001011111110111;
            12'b010111011100: out = 32'b00000000000000111001100011011111;
            12'b010111011101: out = 32'b00000000000000111001100111000110;
            12'b010111011110: out = 32'b00000000000000111001101010101110;
            12'b010111011111: out = 32'b00000000000000111001101110010110;
            12'b010111100000: out = 32'b00000000000000111001110001111110;
            12'b010111100001: out = 32'b00000000000000111001110101100111;
            12'b010111100010: out = 32'b00000000000000111001111001001111;
            12'b010111100011: out = 32'b00000000000000111001111100111000;
            12'b010111100100: out = 32'b00000000000000111010000000100001;
            12'b010111100101: out = 32'b00000000000000111010000100001011;
            12'b010111100110: out = 32'b00000000000000111010000111110100;
            12'b010111100111: out = 32'b00000000000000111010001011011110;
            12'b010111101000: out = 32'b00000000000000111010001111001000;
            12'b010111101001: out = 32'b00000000000000111010010010110010;
            12'b010111101010: out = 32'b00000000000000111010010110011100;
            12'b010111101011: out = 32'b00000000000000111010011010000110;
            12'b010111101100: out = 32'b00000000000000111010011101110001;
            12'b010111101101: out = 32'b00000000000000111010100001011100;
            12'b010111101110: out = 32'b00000000000000111010100101000111;
            12'b010111101111: out = 32'b00000000000000111010101000110011;
            12'b010111110000: out = 32'b00000000000000111010101100011110;
            12'b010111110001: out = 32'b00000000000000111010110000001010;
            12'b010111110010: out = 32'b00000000000000111010110011110110;
            12'b010111110011: out = 32'b00000000000000111010110111100010;
            12'b010111110100: out = 32'b00000000000000111010111011001110;
            12'b010111110101: out = 32'b00000000000000111010111110111011;
            12'b010111110110: out = 32'b00000000000000111011000010101000;
            12'b010111110111: out = 32'b00000000000000111011000110010101;
            12'b010111111000: out = 32'b00000000000000111011001010000010;
            12'b010111111001: out = 32'b00000000000000111011001101110000;
            12'b010111111010: out = 32'b00000000000000111011010001011101;
            12'b010111111011: out = 32'b00000000000000111011010101001011;
            12'b010111111100: out = 32'b00000000000000111011011000111001;
            12'b010111111101: out = 32'b00000000000000111011011100101000;
            12'b010111111110: out = 32'b00000000000000111011100000010110;
            12'b010111111111: out = 32'b00000000000000111011100100000101;
            12'b011000000000: out = 32'b00000000000000111011100111110100;
            12'b011000000001: out = 32'b00000000000000111011101011100011;
            12'b011000000010: out = 32'b00000000000000111011101111010011;
            12'b011000000011: out = 32'b00000000000000111011110011000010;
            12'b011000000100: out = 32'b00000000000000111011110110110010;
            12'b011000000101: out = 32'b00000000000000111011111010100010;
            12'b011000000110: out = 32'b00000000000000111011111110010010;
            12'b011000000111: out = 32'b00000000000000111100000010000011;
            12'b011000001000: out = 32'b00000000000000111100000101110100;
            12'b011000001001: out = 32'b00000000000000111100001001100101;
            12'b011000001010: out = 32'b00000000000000111100001101010110;
            12'b011000001011: out = 32'b00000000000000111100010001000111;
            12'b011000001100: out = 32'b00000000000000111100010100111001;
            12'b011000001101: out = 32'b00000000000000111100011000101011;
            12'b011000001110: out = 32'b00000000000000111100011100011101;
            12'b011000001111: out = 32'b00000000000000111100100000001111;
            12'b011000010000: out = 32'b00000000000000111100100100000001;
            12'b011000010001: out = 32'b00000000000000111100100111110100;
            12'b011000010010: out = 32'b00000000000000111100101011100111;
            12'b011000010011: out = 32'b00000000000000111100101111011010;
            12'b011000010100: out = 32'b00000000000000111100110011001110;
            12'b011000010101: out = 32'b00000000000000111100110111000001;
            12'b011000010110: out = 32'b00000000000000111100111010110101;
            12'b011000010111: out = 32'b00000000000000111100111110101001;
            12'b011000011000: out = 32'b00000000000000111101000010011110;
            12'b011000011001: out = 32'b00000000000000111101000110010010;
            12'b011000011010: out = 32'b00000000000000111101001010000111;
            12'b011000011011: out = 32'b00000000000000111101001101111100;
            12'b011000011100: out = 32'b00000000000000111101010001110001;
            12'b011000011101: out = 32'b00000000000000111101010101100111;
            12'b011000011110: out = 32'b00000000000000111101011001011100;
            12'b011000011111: out = 32'b00000000000000111101011101010010;
            12'b011000100000: out = 32'b00000000000000111101100001001000;
            12'b011000100001: out = 32'b00000000000000111101100100111111;
            12'b011000100010: out = 32'b00000000000000111101101000110101;
            12'b011000100011: out = 32'b00000000000000111101101100101100;
            12'b011000100100: out = 32'b00000000000000111101110000100011;
            12'b011000100101: out = 32'b00000000000000111101110100011011;
            12'b011000100110: out = 32'b00000000000000111101111000010010;
            12'b011000100111: out = 32'b00000000000000111101111100001010;
            12'b011000101000: out = 32'b00000000000000111110000000000010;
            12'b011000101001: out = 32'b00000000000000111110000011111010;
            12'b011000101010: out = 32'b00000000000000111110000111110011;
            12'b011000101011: out = 32'b00000000000000111110001011101011;
            12'b011000101100: out = 32'b00000000000000111110001111100100;
            12'b011000101101: out = 32'b00000000000000111110010011011110;
            12'b011000101110: out = 32'b00000000000000111110010111010111;
            12'b011000101111: out = 32'b00000000000000111110011011010001;
            12'b011000110000: out = 32'b00000000000000111110011111001010;
            12'b011000110001: out = 32'b00000000000000111110100011000101;
            12'b011000110010: out = 32'b00000000000000111110100110111111;
            12'b011000110011: out = 32'b00000000000000111110101010111010;
            12'b011000110100: out = 32'b00000000000000111110101110110100;
            12'b011000110101: out = 32'b00000000000000111110110010110000;
            12'b011000110110: out = 32'b00000000000000111110110110101011;
            12'b011000110111: out = 32'b00000000000000111110111010100110;
            12'b011000111000: out = 32'b00000000000000111110111110100010;
            12'b011000111001: out = 32'b00000000000000111111000010011110;
            12'b011000111010: out = 32'b00000000000000111111000110011011;
            12'b011000111011: out = 32'b00000000000000111111001010010111;
            12'b011000111100: out = 32'b00000000000000111111001110010100;
            12'b011000111101: out = 32'b00000000000000111111010010010001;
            12'b011000111110: out = 32'b00000000000000111111010110001110;
            12'b011000111111: out = 32'b00000000000000111111011010001100;
            12'b011001000000: out = 32'b00000000000000111111011110001010;
            12'b011001000001: out = 32'b00000000000000111111100010001000;
            12'b011001000010: out = 32'b00000000000000111111100110000110;
            12'b011001000011: out = 32'b00000000000000111111101010000100;
            12'b011001000100: out = 32'b00000000000000111111101110000011;
            12'b011001000101: out = 32'b00000000000000111111110010000010;
            12'b011001000110: out = 32'b00000000000000111111110110000001;
            12'b011001000111: out = 32'b00000000000000111111111010000001;
            12'b011001001000: out = 32'b00000000000000111111111110000001;
            default: out = 0;
        endcase
    end
endmodule: tangent_lut
