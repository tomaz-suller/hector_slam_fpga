module cossine_lut
(
    input logic [31:0] in,
    output logic [31:0] out
);

    logic [11:0] truncated_in;
    assign truncated_in = in [18:7];

    always_comb begin
        case (truncated_in)
            12'b000000000000: out = 32'b00000000000001000000000000000000;
            12'b000000000001: out = 32'b00000000000000111111111111111111;
            12'b000000000010: out = 32'b00000000000000111111111111111111;
            12'b000000000011: out = 32'b00000000000000111111111111111111;
            12'b000000000100: out = 32'b00000000000000111111111111111111;
            12'b000000000101: out = 32'b00000000000000111111111111111111;
            12'b000000000110: out = 32'b00000000000000111111111111111110;
            12'b000000000111: out = 32'b00000000000000111111111111111110;
            12'b000000001000: out = 32'b00000000000000111111111111111110;
            12'b000000001001: out = 32'b00000000000000111111111111111101;
            12'b000000001010: out = 32'b00000000000000111111111111111100;
            12'b000000001011: out = 32'b00000000000000111111111111111100;
            12'b000000001100: out = 32'b00000000000000111111111111111011;
            12'b000000001101: out = 32'b00000000000000111111111111111010;
            12'b000000001110: out = 32'b00000000000000111111111111111001;
            12'b000000001111: out = 32'b00000000000000111111111111111000;
            12'b000000010000: out = 32'b00000000000000111111111111111000;
            12'b000000010001: out = 32'b00000000000000111111111111110110;
            12'b000000010010: out = 32'b00000000000000111111111111110101;
            12'b000000010011: out = 32'b00000000000000111111111111110100;
            12'b000000010100: out = 32'b00000000000000111111111111110011;
            12'b000000010101: out = 32'b00000000000000111111111111110010;
            12'b000000010110: out = 32'b00000000000000111111111111110000;
            12'b000000010111: out = 32'b00000000000000111111111111101111;
            12'b000000011000: out = 32'b00000000000000111111111111101110;
            12'b000000011001: out = 32'b00000000000000111111111111101100;
            12'b000000011010: out = 32'b00000000000000111111111111101010;
            12'b000000011011: out = 32'b00000000000000111111111111101001;
            12'b000000011100: out = 32'b00000000000000111111111111100111;
            12'b000000011101: out = 32'b00000000000000111111111111100101;
            12'b000000011110: out = 32'b00000000000000111111111111100011;
            12'b000000011111: out = 32'b00000000000000111111111111100001;
            12'b000000100000: out = 32'b00000000000000111111111111100000;
            12'b000000100001: out = 32'b00000000000000111111111111011101;
            12'b000000100010: out = 32'b00000000000000111111111111011011;
            12'b000000100011: out = 32'b00000000000000111111111111011001;
            12'b000000100100: out = 32'b00000000000000111111111111010111;
            12'b000000100101: out = 32'b00000000000000111111111111010101;
            12'b000000100110: out = 32'b00000000000000111111111111010010;
            12'b000000100111: out = 32'b00000000000000111111111111010000;
            12'b000000101000: out = 32'b00000000000000111111111111001110;
            12'b000000101001: out = 32'b00000000000000111111111111001011;
            12'b000000101010: out = 32'b00000000000000111111111111001000;
            12'b000000101011: out = 32'b00000000000000111111111111000110;
            12'b000000101100: out = 32'b00000000000000111111111111000011;
            12'b000000101101: out = 32'b00000000000000111111111111000000;
            12'b000000101110: out = 32'b00000000000000111111111110111101;
            12'b000000101111: out = 32'b00000000000000111111111110111010;
            12'b000000110000: out = 32'b00000000000000111111111110111000;
            12'b000000110001: out = 32'b00000000000000111111111110110100;
            12'b000000110010: out = 32'b00000000000000111111111110110001;
            12'b000000110011: out = 32'b00000000000000111111111110101110;
            12'b000000110100: out = 32'b00000000000000111111111110101011;
            12'b000000110101: out = 32'b00000000000000111111111110101000;
            12'b000000110110: out = 32'b00000000000000111111111110100100;
            12'b000000110111: out = 32'b00000000000000111111111110100001;
            12'b000000111000: out = 32'b00000000000000111111111110011110;
            12'b000000111001: out = 32'b00000000000000111111111110011010;
            12'b000000111010: out = 32'b00000000000000111111111110010110;
            12'b000000111011: out = 32'b00000000000000111111111110010011;
            12'b000000111100: out = 32'b00000000000000111111111110001111;
            12'b000000111101: out = 32'b00000000000000111111111110001011;
            12'b000000111110: out = 32'b00000000000000111111111110000111;
            12'b000000111111: out = 32'b00000000000000111111111110000011;
            12'b000001000000: out = 32'b00000000000000111111111110000000;
            12'b000001000001: out = 32'b00000000000000111111111101111011;
            12'b000001000010: out = 32'b00000000000000111111111101110111;
            12'b000001000011: out = 32'b00000000000000111111111101110011;
            12'b000001000100: out = 32'b00000000000000111111111101101111;
            12'b000001000101: out = 32'b00000000000000111111111101101011;
            12'b000001000110: out = 32'b00000000000000111111111101100110;
            12'b000001000111: out = 32'b00000000000000111111111101100010;
            12'b000001001000: out = 32'b00000000000000111111111101011110;
            12'b000001001001: out = 32'b00000000000000111111111101011001;
            12'b000001001010: out = 32'b00000000000000111111111101010100;
            12'b000001001011: out = 32'b00000000000000111111111101010000;
            12'b000001001100: out = 32'b00000000000000111111111101001011;
            12'b000001001101: out = 32'b00000000000000111111111101000110;
            12'b000001001110: out = 32'b00000000000000111111111101000001;
            12'b000001001111: out = 32'b00000000000000111111111100111100;
            12'b000001010000: out = 32'b00000000000000111111111100111000;
            12'b000001010001: out = 32'b00000000000000111111111100110010;
            12'b000001010010: out = 32'b00000000000000111111111100101101;
            12'b000001010011: out = 32'b00000000000000111111111100101000;
            12'b000001010100: out = 32'b00000000000000111111111100100011;
            12'b000001010101: out = 32'b00000000000000111111111100011110;
            12'b000001010110: out = 32'b00000000000000111111111100011000;
            12'b000001010111: out = 32'b00000000000000111111111100010011;
            12'b000001011000: out = 32'b00000000000000111111111100001110;
            12'b000001011001: out = 32'b00000000000000111111111100001000;
            12'b000001011010: out = 32'b00000000000000111111111100000010;
            12'b000001011011: out = 32'b00000000000000111111111011111101;
            12'b000001011100: out = 32'b00000000000000111111111011110111;
            12'b000001011101: out = 32'b00000000000000111111111011110001;
            12'b000001011110: out = 32'b00000000000000111111111011101011;
            12'b000001011111: out = 32'b00000000000000111111111011100110;
            12'b000001100000: out = 32'b00000000000000111111111011100000;
            12'b000001100001: out = 32'b00000000000000111111111011011010;
            12'b000001100010: out = 32'b00000000000000111111111011010011;
            12'b000001100011: out = 32'b00000000000000111111111011001101;
            12'b000001100100: out = 32'b00000000000000111111111011000111;
            12'b000001100101: out = 32'b00000000000000111111111011000001;
            12'b000001100110: out = 32'b00000000000000111111111010111010;
            12'b000001100111: out = 32'b00000000000000111111111010110100;
            12'b000001101000: out = 32'b00000000000000111111111010101110;
            12'b000001101001: out = 32'b00000000000000111111111010100111;
            12'b000001101010: out = 32'b00000000000000111111111010100000;
            12'b000001101011: out = 32'b00000000000000111111111010011010;
            12'b000001101100: out = 32'b00000000000000111111111010010011;
            12'b000001101101: out = 32'b00000000000000111111111010001100;
            12'b000001101110: out = 32'b00000000000000111111111010000101;
            12'b000001101111: out = 32'b00000000000000111111111001111111;
            12'b000001110000: out = 32'b00000000000000111111111001111000;
            12'b000001110001: out = 32'b00000000000000111111111001110001;
            12'b000001110010: out = 32'b00000000000000111111111001101001;
            12'b000001110011: out = 32'b00000000000000111111111001100010;
            12'b000001110100: out = 32'b00000000000000111111111001011011;
            12'b000001110101: out = 32'b00000000000000111111111001010100;
            12'b000001110110: out = 32'b00000000000000111111111001001100;
            12'b000001110111: out = 32'b00000000000000111111111001000101;
            12'b000001111000: out = 32'b00000000000000111111111000111110;
            12'b000001111001: out = 32'b00000000000000111111111000110110;
            12'b000001111010: out = 32'b00000000000000111111111000101111;
            12'b000001111011: out = 32'b00000000000000111111111000100111;
            12'b000001111100: out = 32'b00000000000000111111111000011111;
            12'b000001111101: out = 32'b00000000000000111111111000010111;
            12'b000001111110: out = 32'b00000000000000111111111000010000;
            12'b000001111111: out = 32'b00000000000000111111111000001000;
            12'b000010000000: out = 32'b00000000000000111111111000000000;
            12'b000010000001: out = 32'b00000000000000111111110111111000;
            12'b000010000010: out = 32'b00000000000000111111110111110000;
            12'b000010000011: out = 32'b00000000000000111111110111100111;
            12'b000010000100: out = 32'b00000000000000111111110111011111;
            12'b000010000101: out = 32'b00000000000000111111110111010111;
            12'b000010000110: out = 32'b00000000000000111111110111001111;
            12'b000010000111: out = 32'b00000000000000111111110111000110;
            12'b000010001000: out = 32'b00000000000000111111110110111110;
            12'b000010001001: out = 32'b00000000000000111111110110110101;
            12'b000010001010: out = 32'b00000000000000111111110110101101;
            12'b000010001011: out = 32'b00000000000000111111110110100100;
            12'b000010001100: out = 32'b00000000000000111111110110011011;
            12'b000010001101: out = 32'b00000000000000111111110110010010;
            12'b000010001110: out = 32'b00000000000000111111110110001010;
            12'b000010001111: out = 32'b00000000000000111111110110000001;
            12'b000010010000: out = 32'b00000000000000111111110101111000;
            12'b000010010001: out = 32'b00000000000000111111110101101111;
            12'b000010010010: out = 32'b00000000000000111111110101100110;
            12'b000010010011: out = 32'b00000000000000111111110101011101;
            12'b000010010100: out = 32'b00000000000000111111110101010011;
            12'b000010010101: out = 32'b00000000000000111111110101001010;
            12'b000010010110: out = 32'b00000000000000111111110101000001;
            12'b000010010111: out = 32'b00000000000000111111110100110111;
            12'b000010011000: out = 32'b00000000000000111111110100101110;
            12'b000010011001: out = 32'b00000000000000111111110100100100;
            12'b000010011010: out = 32'b00000000000000111111110100011011;
            12'b000010011011: out = 32'b00000000000000111111110100010001;
            12'b000010011100: out = 32'b00000000000000111111110100000111;
            12'b000010011101: out = 32'b00000000000000111111110011111110;
            12'b000010011110: out = 32'b00000000000000111111110011110100;
            12'b000010011111: out = 32'b00000000000000111111110011101010;
            12'b000010100000: out = 32'b00000000000000111111110011100000;
            12'b000010100001: out = 32'b00000000000000111111110011010110;
            12'b000010100010: out = 32'b00000000000000111111110011001100;
            12'b000010100011: out = 32'b00000000000000111111110011000010;
            12'b000010100100: out = 32'b00000000000000111111110010110111;
            12'b000010100101: out = 32'b00000000000000111111110010101101;
            12'b000010100110: out = 32'b00000000000000111111110010100011;
            12'b000010100111: out = 32'b00000000000000111111110010011000;
            12'b000010101000: out = 32'b00000000000000111111110010001110;
            12'b000010101001: out = 32'b00000000000000111111110010000011;
            12'b000010101010: out = 32'b00000000000000111111110001111001;
            12'b000010101011: out = 32'b00000000000000111111110001101110;
            12'b000010101100: out = 32'b00000000000000111111110001100100;
            12'b000010101101: out = 32'b00000000000000111111110001011001;
            12'b000010101110: out = 32'b00000000000000111111110001001110;
            12'b000010101111: out = 32'b00000000000000111111110001000011;
            12'b000010110000: out = 32'b00000000000000111111110000111000;
            12'b000010110001: out = 32'b00000000000000111111110000101101;
            12'b000010110010: out = 32'b00000000000000111111110000100010;
            12'b000010110011: out = 32'b00000000000000111111110000010111;
            12'b000010110100: out = 32'b00000000000000111111110000001100;
            12'b000010110101: out = 32'b00000000000000111111110000000000;
            12'b000010110110: out = 32'b00000000000000111111101111110101;
            12'b000010110111: out = 32'b00000000000000111111101111101010;
            12'b000010111000: out = 32'b00000000000000111111101111011110;
            12'b000010111001: out = 32'b00000000000000111111101111010011;
            12'b000010111010: out = 32'b00000000000000111111101111000111;
            12'b000010111011: out = 32'b00000000000000111111101110111011;
            12'b000010111100: out = 32'b00000000000000111111101110110000;
            12'b000010111101: out = 32'b00000000000000111111101110100100;
            12'b000010111110: out = 32'b00000000000000111111101110011000;
            12'b000010111111: out = 32'b00000000000000111111101110001100;
            12'b000011000000: out = 32'b00000000000000111111101110000000;
            12'b000011000001: out = 32'b00000000000000111111101101110100;
            12'b000011000010: out = 32'b00000000000000111111101101101000;
            12'b000011000011: out = 32'b00000000000000111111101101011100;
            12'b000011000100: out = 32'b00000000000000111111101101010000;
            12'b000011000101: out = 32'b00000000000000111111101101000100;
            12'b000011000110: out = 32'b00000000000000111111101100110111;
            12'b000011000111: out = 32'b00000000000000111111101100101011;
            12'b000011001000: out = 32'b00000000000000111111101100011110;
            12'b000011001001: out = 32'b00000000000000111111101100010010;
            12'b000011001010: out = 32'b00000000000000111111101100000101;
            12'b000011001011: out = 32'b00000000000000111111101011111001;
            12'b000011001100: out = 32'b00000000000000111111101011101100;
            12'b000011001101: out = 32'b00000000000000111111101011011111;
            12'b000011001110: out = 32'b00000000000000111111101011010010;
            12'b000011001111: out = 32'b00000000000000111111101011000110;
            12'b000011010000: out = 32'b00000000000000111111101010111001;
            12'b000011010001: out = 32'b00000000000000111111101010101100;
            12'b000011010010: out = 32'b00000000000000111111101010011111;
            12'b000011010011: out = 32'b00000000000000111111101010010001;
            12'b000011010100: out = 32'b00000000000000111111101010000100;
            12'b000011010101: out = 32'b00000000000000111111101001110111;
            12'b000011010110: out = 32'b00000000000000111111101001101010;
            12'b000011010111: out = 32'b00000000000000111111101001011100;
            12'b000011011000: out = 32'b00000000000000111111101001001111;
            12'b000011011001: out = 32'b00000000000000111111101001000001;
            12'b000011011010: out = 32'b00000000000000111111101000110100;
            12'b000011011011: out = 32'b00000000000000111111101000100110;
            12'b000011011100: out = 32'b00000000000000111111101000011000;
            12'b000011011101: out = 32'b00000000000000111111101000001011;
            12'b000011011110: out = 32'b00000000000000111111100111111101;
            12'b000011011111: out = 32'b00000000000000111111100111101111;
            12'b000011100000: out = 32'b00000000000000111111100111100001;
            12'b000011100001: out = 32'b00000000000000111111100111010011;
            12'b000011100010: out = 32'b00000000000000111111100111000101;
            12'b000011100011: out = 32'b00000000000000111111100110110111;
            12'b000011100100: out = 32'b00000000000000111111100110101001;
            12'b000011100101: out = 32'b00000000000000111111100110011010;
            12'b000011100110: out = 32'b00000000000000111111100110001100;
            12'b000011100111: out = 32'b00000000000000111111100101111110;
            12'b000011101000: out = 32'b00000000000000111111100101101111;
            12'b000011101001: out = 32'b00000000000000111111100101100001;
            12'b000011101010: out = 32'b00000000000000111111100101010010;
            12'b000011101011: out = 32'b00000000000000111111100101000100;
            12'b000011101100: out = 32'b00000000000000111111100100110101;
            12'b000011101101: out = 32'b00000000000000111111100100100110;
            12'b000011101110: out = 32'b00000000000000111111100100010111;
            12'b000011101111: out = 32'b00000000000000111111100100001000;
            12'b000011110000: out = 32'b00000000000000111111100011111010;
            12'b000011110001: out = 32'b00000000000000111111100011101011;
            12'b000011110010: out = 32'b00000000000000111111100011011100;
            12'b000011110011: out = 32'b00000000000000111111100011001100;
            12'b000011110100: out = 32'b00000000000000111111100010111101;
            12'b000011110101: out = 32'b00000000000000111111100010101110;
            12'b000011110110: out = 32'b00000000000000111111100010011111;
            12'b000011110111: out = 32'b00000000000000111111100010001111;
            12'b000011111000: out = 32'b00000000000000111111100010000000;
            12'b000011111001: out = 32'b00000000000000111111100001110000;
            12'b000011111010: out = 32'b00000000000000111111100001100001;
            12'b000011111011: out = 32'b00000000000000111111100001010001;
            12'b000011111100: out = 32'b00000000000000111111100001000010;
            12'b000011111101: out = 32'b00000000000000111111100000110010;
            12'b000011111110: out = 32'b00000000000000111111100000100010;
            12'b000011111111: out = 32'b00000000000000111111100000010010;
            12'b000100000000: out = 32'b00000000000000111111100000000010;
            12'b000100000001: out = 32'b00000000000000111111011111110010;
            12'b000100000010: out = 32'b00000000000000111111011111100010;
            12'b000100000011: out = 32'b00000000000000111111011111010010;
            12'b000100000100: out = 32'b00000000000000111111011111000010;
            12'b000100000101: out = 32'b00000000000000111111011110110010;
            12'b000100000110: out = 32'b00000000000000111111011110100001;
            12'b000100000111: out = 32'b00000000000000111111011110010001;
            12'b000100001000: out = 32'b00000000000000111111011110000001;
            12'b000100001001: out = 32'b00000000000000111111011101110000;
            12'b000100001010: out = 32'b00000000000000111111011101011111;
            12'b000100001011: out = 32'b00000000000000111111011101001111;
            12'b000100001100: out = 32'b00000000000000111111011100111110;
            12'b000100001101: out = 32'b00000000000000111111011100101101;
            12'b000100001110: out = 32'b00000000000000111111011100011101;
            12'b000100001111: out = 32'b00000000000000111111011100001100;
            12'b000100010000: out = 32'b00000000000000111111011011111011;
            12'b000100010001: out = 32'b00000000000000111111011011101010;
            12'b000100010010: out = 32'b00000000000000111111011011011001;
            12'b000100010011: out = 32'b00000000000000111111011011001000;
            12'b000100010100: out = 32'b00000000000000111111011010110111;
            12'b000100010101: out = 32'b00000000000000111111011010100101;
            12'b000100010110: out = 32'b00000000000000111111011010010100;
            12'b000100010111: out = 32'b00000000000000111111011010000011;
            12'b000100011000: out = 32'b00000000000000111111011001110001;
            12'b000100011001: out = 32'b00000000000000111111011001100000;
            12'b000100011010: out = 32'b00000000000000111111011001001110;
            12'b000100011011: out = 32'b00000000000000111111011000111101;
            12'b000100011100: out = 32'b00000000000000111111011000101011;
            12'b000100011101: out = 32'b00000000000000111111011000011001;
            12'b000100011110: out = 32'b00000000000000111111011000001000;
            12'b000100011111: out = 32'b00000000000000111111010111110110;
            12'b000100100000: out = 32'b00000000000000111111010111100100;
            12'b000100100001: out = 32'b00000000000000111111010111010010;
            12'b000100100010: out = 32'b00000000000000111111010111000000;
            12'b000100100011: out = 32'b00000000000000111111010110101110;
            12'b000100100100: out = 32'b00000000000000111111010110011100;
            12'b000100100101: out = 32'b00000000000000111111010110001001;
            12'b000100100110: out = 32'b00000000000000111111010101110111;
            12'b000100100111: out = 32'b00000000000000111111010101100101;
            12'b000100101000: out = 32'b00000000000000111111010101010010;
            12'b000100101001: out = 32'b00000000000000111111010101000000;
            12'b000100101010: out = 32'b00000000000000111111010100101101;
            12'b000100101011: out = 32'b00000000000000111111010100011011;
            12'b000100101100: out = 32'b00000000000000111111010100001000;
            12'b000100101101: out = 32'b00000000000000111111010011110101;
            12'b000100101110: out = 32'b00000000000000111111010011100011;
            12'b000100101111: out = 32'b00000000000000111111010011010000;
            12'b000100110000: out = 32'b00000000000000111111010010111101;
            12'b000100110001: out = 32'b00000000000000111111010010101010;
            12'b000100110010: out = 32'b00000000000000111111010010010111;
            12'b000100110011: out = 32'b00000000000000111111010010000100;
            12'b000100110100: out = 32'b00000000000000111111010001110001;
            12'b000100110101: out = 32'b00000000000000111111010001011101;
            12'b000100110110: out = 32'b00000000000000111111010001001010;
            12'b000100110111: out = 32'b00000000000000111111010000110111;
            12'b000100111000: out = 32'b00000000000000111111010000100011;
            12'b000100111001: out = 32'b00000000000000111111010000010000;
            12'b000100111010: out = 32'b00000000000000111111001111111100;
            12'b000100111011: out = 32'b00000000000000111111001111101001;
            12'b000100111100: out = 32'b00000000000000111111001111010101;
            12'b000100111101: out = 32'b00000000000000111111001111000001;
            12'b000100111110: out = 32'b00000000000000111111001110101110;
            12'b000100111111: out = 32'b00000000000000111111001110011010;
            12'b000101000000: out = 32'b00000000000000111111001110000110;
            12'b000101000001: out = 32'b00000000000000111111001101110010;
            12'b000101000010: out = 32'b00000000000000111111001101011110;
            12'b000101000011: out = 32'b00000000000000111111001101001010;
            12'b000101000100: out = 32'b00000000000000111111001100110110;
            12'b000101000101: out = 32'b00000000000000111111001100100010;
            12'b000101000110: out = 32'b00000000000000111111001100001101;
            12'b000101000111: out = 32'b00000000000000111111001011111001;
            12'b000101001000: out = 32'b00000000000000111111001011100101;
            12'b000101001001: out = 32'b00000000000000111111001011010000;
            12'b000101001010: out = 32'b00000000000000111111001010111100;
            12'b000101001011: out = 32'b00000000000000111111001010100111;
            12'b000101001100: out = 32'b00000000000000111111001010010011;
            12'b000101001101: out = 32'b00000000000000111111001001111110;
            12'b000101001110: out = 32'b00000000000000111111001001101001;
            12'b000101001111: out = 32'b00000000000000111111001001010100;
            12'b000101010000: out = 32'b00000000000000111111001000111111;
            12'b000101010001: out = 32'b00000000000000111111001000101010;
            12'b000101010010: out = 32'b00000000000000111111001000010101;
            12'b000101010011: out = 32'b00000000000000111111001000000000;
            12'b000101010100: out = 32'b00000000000000111111000111101011;
            12'b000101010101: out = 32'b00000000000000111111000111010110;
            12'b000101010110: out = 32'b00000000000000111111000111000001;
            12'b000101010111: out = 32'b00000000000000111111000110101100;
            12'b000101011000: out = 32'b00000000000000111111000110010110;
            12'b000101011001: out = 32'b00000000000000111111000110000001;
            12'b000101011010: out = 32'b00000000000000111111000101101011;
            12'b000101011011: out = 32'b00000000000000111111000101010110;
            12'b000101011100: out = 32'b00000000000000111111000101000000;
            12'b000101011101: out = 32'b00000000000000111111000100101010;
            12'b000101011110: out = 32'b00000000000000111111000100010101;
            12'b000101011111: out = 32'b00000000000000111111000011111111;
            12'b000101100000: out = 32'b00000000000000111111000011101001;
            12'b000101100001: out = 32'b00000000000000111111000011010011;
            12'b000101100010: out = 32'b00000000000000111111000010111101;
            12'b000101100011: out = 32'b00000000000000111111000010100111;
            12'b000101100100: out = 32'b00000000000000111111000010010001;
            12'b000101100101: out = 32'b00000000000000111111000001111011;
            12'b000101100110: out = 32'b00000000000000111111000001100101;
            12'b000101100111: out = 32'b00000000000000111111000001001110;
            12'b000101101000: out = 32'b00000000000000111111000000111000;
            12'b000101101001: out = 32'b00000000000000111111000000100010;
            12'b000101101010: out = 32'b00000000000000111111000000001011;
            12'b000101101011: out = 32'b00000000000000111110111111110100;
            12'b000101101100: out = 32'b00000000000000111110111111011110;
            12'b000101101101: out = 32'b00000000000000111110111111000111;
            12'b000101101110: out = 32'b00000000000000111110111110110001;
            12'b000101101111: out = 32'b00000000000000111110111110011010;
            12'b000101110000: out = 32'b00000000000000111110111110000011;
            12'b000101110001: out = 32'b00000000000000111110111101101100;
            12'b000101110010: out = 32'b00000000000000111110111101010101;
            12'b000101110011: out = 32'b00000000000000111110111100111110;
            12'b000101110100: out = 32'b00000000000000111110111100100111;
            12'b000101110101: out = 32'b00000000000000111110111100010000;
            12'b000101110110: out = 32'b00000000000000111110111011111001;
            12'b000101110111: out = 32'b00000000000000111110111011100001;
            12'b000101111000: out = 32'b00000000000000111110111011001010;
            12'b000101111001: out = 32'b00000000000000111110111010110010;
            12'b000101111010: out = 32'b00000000000000111110111010011011;
            12'b000101111011: out = 32'b00000000000000111110111010000100;
            12'b000101111100: out = 32'b00000000000000111110111001101100;
            12'b000101111101: out = 32'b00000000000000111110111001010100;
            12'b000101111110: out = 32'b00000000000000111110111000111101;
            12'b000101111111: out = 32'b00000000000000111110111000100101;
            12'b000110000000: out = 32'b00000000000000111110111000001101;
            12'b000110000001: out = 32'b00000000000000111110110111110101;
            12'b000110000010: out = 32'b00000000000000111110110111011101;
            12'b000110000011: out = 32'b00000000000000111110110111000101;
            12'b000110000100: out = 32'b00000000000000111110110110101101;
            12'b000110000101: out = 32'b00000000000000111110110110010101;
            12'b000110000110: out = 32'b00000000000000111110110101111101;
            12'b000110000111: out = 32'b00000000000000111110110101100100;
            12'b000110001000: out = 32'b00000000000000111110110101001100;
            12'b000110001001: out = 32'b00000000000000111110110100110100;
            12'b000110001010: out = 32'b00000000000000111110110100011011;
            12'b000110001011: out = 32'b00000000000000111110110100000011;
            12'b000110001100: out = 32'b00000000000000111110110011101010;
            12'b000110001101: out = 32'b00000000000000111110110011010010;
            12'b000110001110: out = 32'b00000000000000111110110010111001;
            12'b000110001111: out = 32'b00000000000000111110110010100000;
            12'b000110010000: out = 32'b00000000000000111110110010000111;
            12'b000110010001: out = 32'b00000000000000111110110001101111;
            12'b000110010010: out = 32'b00000000000000111110110001010110;
            12'b000110010011: out = 32'b00000000000000111110110000111101;
            12'b000110010100: out = 32'b00000000000000111110110000100100;
            12'b000110010101: out = 32'b00000000000000111110110000001010;
            12'b000110010110: out = 32'b00000000000000111110101111110001;
            12'b000110010111: out = 32'b00000000000000111110101111011000;
            12'b000110011000: out = 32'b00000000000000111110101110111111;
            12'b000110011001: out = 32'b00000000000000111110101110100101;
            12'b000110011010: out = 32'b00000000000000111110101110001100;
            12'b000110011011: out = 32'b00000000000000111110101101110010;
            12'b000110011100: out = 32'b00000000000000111110101101011001;
            12'b000110011101: out = 32'b00000000000000111110101100111111;
            12'b000110011110: out = 32'b00000000000000111110101100100110;
            12'b000110011111: out = 32'b00000000000000111110101100001100;
            12'b000110100000: out = 32'b00000000000000111110101011110010;
            12'b000110100001: out = 32'b00000000000000111110101011011000;
            12'b000110100010: out = 32'b00000000000000111110101010111110;
            12'b000110100011: out = 32'b00000000000000111110101010100100;
            12'b000110100100: out = 32'b00000000000000111110101010001010;
            12'b000110100101: out = 32'b00000000000000111110101001110000;
            12'b000110100110: out = 32'b00000000000000111110101001010110;
            12'b000110100111: out = 32'b00000000000000111110101000111100;
            12'b000110101000: out = 32'b00000000000000111110101000100010;
            12'b000110101001: out = 32'b00000000000000111110101000000111;
            12'b000110101010: out = 32'b00000000000000111110100111101101;
            12'b000110101011: out = 32'b00000000000000111110100111010010;
            12'b000110101100: out = 32'b00000000000000111110100110111000;
            12'b000110101101: out = 32'b00000000000000111110100110011101;
            12'b000110101110: out = 32'b00000000000000111110100110000011;
            12'b000110101111: out = 32'b00000000000000111110100101101000;
            12'b000110110000: out = 32'b00000000000000111110100101001101;
            12'b000110110001: out = 32'b00000000000000111110100100110010;
            12'b000110110010: out = 32'b00000000000000111110100100010111;
            12'b000110110011: out = 32'b00000000000000111110100011111100;
            12'b000110110100: out = 32'b00000000000000111110100011100001;
            12'b000110110101: out = 32'b00000000000000111110100011000110;
            12'b000110110110: out = 32'b00000000000000111110100010101011;
            12'b000110110111: out = 32'b00000000000000111110100010010000;
            12'b000110111000: out = 32'b00000000000000111110100001110101;
            12'b000110111001: out = 32'b00000000000000111110100001011001;
            12'b000110111010: out = 32'b00000000000000111110100000111110;
            12'b000110111011: out = 32'b00000000000000111110100000100011;
            12'b000110111100: out = 32'b00000000000000111110100000000111;
            12'b000110111101: out = 32'b00000000000000111110011111101100;
            12'b000110111110: out = 32'b00000000000000111110011111010000;
            12'b000110111111: out = 32'b00000000000000111110011110110100;
            12'b000111000000: out = 32'b00000000000000111110011110011000;
            12'b000111000001: out = 32'b00000000000000111110011101111101;
            12'b000111000010: out = 32'b00000000000000111110011101100001;
            12'b000111000011: out = 32'b00000000000000111110011101000101;
            12'b000111000100: out = 32'b00000000000000111110011100101001;
            12'b000111000101: out = 32'b00000000000000111110011100001101;
            12'b000111000110: out = 32'b00000000000000111110011011110001;
            12'b000111000111: out = 32'b00000000000000111110011011010101;
            12'b000111001000: out = 32'b00000000000000111110011010111000;
            12'b000111001001: out = 32'b00000000000000111110011010011100;
            12'b000111001010: out = 32'b00000000000000111110011010000000;
            12'b000111001011: out = 32'b00000000000000111110011001100011;
            12'b000111001100: out = 32'b00000000000000111110011001000111;
            12'b000111001101: out = 32'b00000000000000111110011000101010;
            12'b000111001110: out = 32'b00000000000000111110011000001110;
            12'b000111001111: out = 32'b00000000000000111110010111110001;
            12'b000111010000: out = 32'b00000000000000111110010111010100;
            12'b000111010001: out = 32'b00000000000000111110010110110111;
            12'b000111010010: out = 32'b00000000000000111110010110011011;
            12'b000111010011: out = 32'b00000000000000111110010101111110;
            12'b000111010100: out = 32'b00000000000000111110010101100001;
            12'b000111010101: out = 32'b00000000000000111110010101000100;
            12'b000111010110: out = 32'b00000000000000111110010100100111;
            12'b000111010111: out = 32'b00000000000000111110010100001001;
            12'b000111011000: out = 32'b00000000000000111110010011101100;
            12'b000111011001: out = 32'b00000000000000111110010011001111;
            12'b000111011010: out = 32'b00000000000000111110010010110010;
            12'b000111011011: out = 32'b00000000000000111110010010010100;
            12'b000111011100: out = 32'b00000000000000111110010001110111;
            12'b000111011101: out = 32'b00000000000000111110010001011001;
            12'b000111011110: out = 32'b00000000000000111110010000111100;
            12'b000111011111: out = 32'b00000000000000111110010000011110;
            12'b000111100000: out = 32'b00000000000000111110010000000000;
            12'b000111100001: out = 32'b00000000000000111110001111100011;
            12'b000111100010: out = 32'b00000000000000111110001111000101;
            12'b000111100011: out = 32'b00000000000000111110001110100111;
            12'b000111100100: out = 32'b00000000000000111110001110001001;
            12'b000111100101: out = 32'b00000000000000111110001101101011;
            12'b000111100110: out = 32'b00000000000000111110001101001101;
            12'b000111100111: out = 32'b00000000000000111110001100101111;
            12'b000111101000: out = 32'b00000000000000111110001100010001;
            12'b000111101001: out = 32'b00000000000000111110001011110010;
            12'b000111101010: out = 32'b00000000000000111110001011010100;
            12'b000111101011: out = 32'b00000000000000111110001010110110;
            12'b000111101100: out = 32'b00000000000000111110001010010111;
            12'b000111101101: out = 32'b00000000000000111110001001111001;
            12'b000111101110: out = 32'b00000000000000111110001001011010;
            12'b000111101111: out = 32'b00000000000000111110001000111100;
            12'b000111110000: out = 32'b00000000000000111110001000011101;
            12'b000111110001: out = 32'b00000000000000111110000111111110;
            12'b000111110010: out = 32'b00000000000000111110000111011111;
            12'b000111110011: out = 32'b00000000000000111110000111000001;
            12'b000111110100: out = 32'b00000000000000111110000110100010;
            12'b000111110101: out = 32'b00000000000000111110000110000011;
            12'b000111110110: out = 32'b00000000000000111110000101100100;
            12'b000111110111: out = 32'b00000000000000111110000101000101;
            12'b000111111000: out = 32'b00000000000000111110000100100101;
            12'b000111111001: out = 32'b00000000000000111110000100000110;
            12'b000111111010: out = 32'b00000000000000111110000011100111;
            12'b000111111011: out = 32'b00000000000000111110000011001000;
            12'b000111111100: out = 32'b00000000000000111110000010101000;
            12'b000111111101: out = 32'b00000000000000111110000010001001;
            12'b000111111110: out = 32'b00000000000000111110000001101001;
            12'b000111111111: out = 32'b00000000000000111110000001001010;
            12'b001000000000: out = 32'b00000000000000111110000000101010;
            12'b001000000001: out = 32'b00000000000000111110000000001010;
            12'b001000000010: out = 32'b00000000000000111101111111101011;
            12'b001000000011: out = 32'b00000000000000111101111111001011;
            12'b001000000100: out = 32'b00000000000000111101111110101011;
            12'b001000000101: out = 32'b00000000000000111101111110001011;
            12'b001000000110: out = 32'b00000000000000111101111101101011;
            12'b001000000111: out = 32'b00000000000000111101111101001011;
            12'b001000001000: out = 32'b00000000000000111101111100101011;
            12'b001000001001: out = 32'b00000000000000111101111100001011;
            12'b001000001010: out = 32'b00000000000000111101111011101010;
            12'b001000001011: out = 32'b00000000000000111101111011001010;
            12'b001000001100: out = 32'b00000000000000111101111010101010;
            12'b001000001101: out = 32'b00000000000000111101111010001001;
            12'b001000001110: out = 32'b00000000000000111101111001101001;
            12'b001000001111: out = 32'b00000000000000111101111001001000;
            12'b001000010000: out = 32'b00000000000000111101111000101000;
            12'b001000010001: out = 32'b00000000000000111101111000000111;
            12'b001000010010: out = 32'b00000000000000111101110111100110;
            12'b001000010011: out = 32'b00000000000000111101110111000101;
            12'b001000010100: out = 32'b00000000000000111101110110100101;
            12'b001000010101: out = 32'b00000000000000111101110110000100;
            12'b001000010110: out = 32'b00000000000000111101110101100011;
            12'b001000010111: out = 32'b00000000000000111101110101000010;
            12'b001000011000: out = 32'b00000000000000111101110100100001;
            12'b001000011001: out = 32'b00000000000000111101110011111111;
            12'b001000011010: out = 32'b00000000000000111101110011011110;
            12'b001000011011: out = 32'b00000000000000111101110010111101;
            12'b001000011100: out = 32'b00000000000000111101110010011100;
            12'b001000011101: out = 32'b00000000000000111101110001111010;
            12'b001000011110: out = 32'b00000000000000111101110001011001;
            12'b001000011111: out = 32'b00000000000000111101110000110111;
            12'b001000100000: out = 32'b00000000000000111101110000010110;
            12'b001000100001: out = 32'b00000000000000111101101111110100;
            12'b001000100010: out = 32'b00000000000000111101101111010010;
            12'b001000100011: out = 32'b00000000000000111101101110110001;
            12'b001000100100: out = 32'b00000000000000111101101110001111;
            12'b001000100101: out = 32'b00000000000000111101101101101101;
            12'b001000100110: out = 32'b00000000000000111101101101001011;
            12'b001000100111: out = 32'b00000000000000111101101100101001;
            12'b001000101000: out = 32'b00000000000000111101101100000111;
            12'b001000101001: out = 32'b00000000000000111101101011100101;
            12'b001000101010: out = 32'b00000000000000111101101011000011;
            12'b001000101011: out = 32'b00000000000000111101101010100000;
            12'b001000101100: out = 32'b00000000000000111101101001111110;
            12'b001000101101: out = 32'b00000000000000111101101001011100;
            12'b001000101110: out = 32'b00000000000000111101101000111001;
            12'b001000101111: out = 32'b00000000000000111101101000010111;
            12'b001000110000: out = 32'b00000000000000111101100111110100;
            12'b001000110001: out = 32'b00000000000000111101100111010010;
            12'b001000110010: out = 32'b00000000000000111101100110101111;
            12'b001000110011: out = 32'b00000000000000111101100110001100;
            12'b001000110100: out = 32'b00000000000000111101100101101010;
            12'b001000110101: out = 32'b00000000000000111101100101000111;
            12'b001000110110: out = 32'b00000000000000111101100100100100;
            12'b001000110111: out = 32'b00000000000000111101100100000001;
            12'b001000111000: out = 32'b00000000000000111101100011011110;
            12'b001000111001: out = 32'b00000000000000111101100010111011;
            12'b001000111010: out = 32'b00000000000000111101100010011000;
            12'b001000111011: out = 32'b00000000000000111101100001110101;
            12'b001000111100: out = 32'b00000000000000111101100001010001;
            12'b001000111101: out = 32'b00000000000000111101100000101110;
            12'b001000111110: out = 32'b00000000000000111101100000001011;
            12'b001000111111: out = 32'b00000000000000111101011111100111;
            12'b001001000000: out = 32'b00000000000000111101011111000100;
            12'b001001000001: out = 32'b00000000000000111101011110100000;
            12'b001001000010: out = 32'b00000000000000111101011101111100;
            12'b001001000011: out = 32'b00000000000000111101011101011001;
            12'b001001000100: out = 32'b00000000000000111101011100110101;
            12'b001001000101: out = 32'b00000000000000111101011100010001;
            12'b001001000110: out = 32'b00000000000000111101011011101101;
            12'b001001000111: out = 32'b00000000000000111101011011001010;
            12'b001001001000: out = 32'b00000000000000111101011010100110;
            12'b001001001001: out = 32'b00000000000000111101011010000001;
            12'b001001001010: out = 32'b00000000000000111101011001011101;
            12'b001001001011: out = 32'b00000000000000111101011000111001;
            12'b001001001100: out = 32'b00000000000000111101011000010101;
            12'b001001001101: out = 32'b00000000000000111101010111110001;
            12'b001001001110: out = 32'b00000000000000111101010111001100;
            12'b001001001111: out = 32'b00000000000000111101010110101000;
            12'b001001010000: out = 32'b00000000000000111101010110000100;
            12'b001001010001: out = 32'b00000000000000111101010101011111;
            12'b001001010010: out = 32'b00000000000000111101010100111010;
            12'b001001010011: out = 32'b00000000000000111101010100010110;
            12'b001001010100: out = 32'b00000000000000111101010011110001;
            12'b001001010101: out = 32'b00000000000000111101010011001100;
            12'b001001010110: out = 32'b00000000000000111101010010101000;
            12'b001001010111: out = 32'b00000000000000111101010010000011;
            12'b001001011000: out = 32'b00000000000000111101010001011110;
            12'b001001011001: out = 32'b00000000000000111101010000111001;
            12'b001001011010: out = 32'b00000000000000111101010000010100;
            12'b001001011011: out = 32'b00000000000000111101001111101111;
            12'b001001011100: out = 32'b00000000000000111101001111001001;
            12'b001001011101: out = 32'b00000000000000111101001110100100;
            12'b001001011110: out = 32'b00000000000000111101001101111111;
            12'b001001011111: out = 32'b00000000000000111101001101011010;
            12'b001001100000: out = 32'b00000000000000111101001100110100;
            12'b001001100001: out = 32'b00000000000000111101001100001111;
            12'b001001100010: out = 32'b00000000000000111101001011101001;
            12'b001001100011: out = 32'b00000000000000111101001011000011;
            12'b001001100100: out = 32'b00000000000000111101001010011110;
            12'b001001100101: out = 32'b00000000000000111101001001111000;
            12'b001001100110: out = 32'b00000000000000111101001001010010;
            12'b001001100111: out = 32'b00000000000000111101001000101101;
            12'b001001101000: out = 32'b00000000000000111101001000000111;
            12'b001001101001: out = 32'b00000000000000111101000111100001;
            12'b001001101010: out = 32'b00000000000000111101000110111011;
            12'b001001101011: out = 32'b00000000000000111101000110010101;
            12'b001001101100: out = 32'b00000000000000111101000101101110;
            12'b001001101101: out = 32'b00000000000000111101000101001000;
            12'b001001101110: out = 32'b00000000000000111101000100100010;
            12'b001001101111: out = 32'b00000000000000111101000011111100;
            12'b001001110000: out = 32'b00000000000000111101000011010101;
            12'b001001110001: out = 32'b00000000000000111101000010101111;
            12'b001001110010: out = 32'b00000000000000111101000010001000;
            12'b001001110011: out = 32'b00000000000000111101000001100010;
            12'b001001110100: out = 32'b00000000000000111101000000111011;
            12'b001001110101: out = 32'b00000000000000111101000000010101;
            12'b001001110110: out = 32'b00000000000000111100111111101110;
            12'b001001110111: out = 32'b00000000000000111100111111000111;
            12'b001001111000: out = 32'b00000000000000111100111110100000;
            12'b001001111001: out = 32'b00000000000000111100111101111001;
            12'b001001111010: out = 32'b00000000000000111100111101010010;
            12'b001001111011: out = 32'b00000000000000111100111100101011;
            12'b001001111100: out = 32'b00000000000000111100111100000100;
            12'b001001111101: out = 32'b00000000000000111100111011011101;
            12'b001001111110: out = 32'b00000000000000111100111010110110;
            12'b001001111111: out = 32'b00000000000000111100111010001111;
            12'b001010000000: out = 32'b00000000000000111100111001100111;
            12'b001010000001: out = 32'b00000000000000111100111001000000;
            12'b001010000010: out = 32'b00000000000000111100111000011001;
            12'b001010000011: out = 32'b00000000000000111100110111110001;
            12'b001010000100: out = 32'b00000000000000111100110111001001;
            12'b001010000101: out = 32'b00000000000000111100110110100010;
            12'b001010000110: out = 32'b00000000000000111100110101111010;
            12'b001010000111: out = 32'b00000000000000111100110101010010;
            12'b001010001000: out = 32'b00000000000000111100110100101011;
            12'b001010001001: out = 32'b00000000000000111100110100000011;
            12'b001010001010: out = 32'b00000000000000111100110011011011;
            12'b001010001011: out = 32'b00000000000000111100110010110011;
            12'b001010001100: out = 32'b00000000000000111100110010001011;
            12'b001010001101: out = 32'b00000000000000111100110001100011;
            12'b001010001110: out = 32'b00000000000000111100110000111011;
            12'b001010001111: out = 32'b00000000000000111100110000010010;
            12'b001010010000: out = 32'b00000000000000111100101111101010;
            12'b001010010001: out = 32'b00000000000000111100101111000010;
            12'b001010010010: out = 32'b00000000000000111100101110011001;
            12'b001010010011: out = 32'b00000000000000111100101101110001;
            12'b001010010100: out = 32'b00000000000000111100101101001000;
            12'b001010010101: out = 32'b00000000000000111100101100100000;
            12'b001010010110: out = 32'b00000000000000111100101011110111;
            12'b001010010111: out = 32'b00000000000000111100101011001111;
            12'b001010011000: out = 32'b00000000000000111100101010100110;
            12'b001010011001: out = 32'b00000000000000111100101001111101;
            12'b001010011010: out = 32'b00000000000000111100101001010100;
            12'b001010011011: out = 32'b00000000000000111100101000101011;
            12'b001010011100: out = 32'b00000000000000111100101000000010;
            12'b001010011101: out = 32'b00000000000000111100100111011001;
            12'b001010011110: out = 32'b00000000000000111100100110110000;
            12'b001010011111: out = 32'b00000000000000111100100110000111;
            12'b001010100000: out = 32'b00000000000000111100100101011110;
            12'b001010100001: out = 32'b00000000000000111100100100110100;
            12'b001010100010: out = 32'b00000000000000111100100100001011;
            12'b001010100011: out = 32'b00000000000000111100100011100010;
            12'b001010100100: out = 32'b00000000000000111100100010111000;
            12'b001010100101: out = 32'b00000000000000111100100010001111;
            12'b001010100110: out = 32'b00000000000000111100100001100101;
            12'b001010100111: out = 32'b00000000000000111100100000111011;
            12'b001010101000: out = 32'b00000000000000111100100000010010;
            12'b001010101001: out = 32'b00000000000000111100011111101000;
            12'b001010101010: out = 32'b00000000000000111100011110111110;
            12'b001010101011: out = 32'b00000000000000111100011110010100;
            12'b001010101100: out = 32'b00000000000000111100011101101010;
            12'b001010101101: out = 32'b00000000000000111100011101000000;
            12'b001010101110: out = 32'b00000000000000111100011100010110;
            12'b001010101111: out = 32'b00000000000000111100011011101100;
            12'b001010110000: out = 32'b00000000000000111100011011000010;
            12'b001010110001: out = 32'b00000000000000111100011010011000;
            12'b001010110010: out = 32'b00000000000000111100011001101110;
            12'b001010110011: out = 32'b00000000000000111100011001000011;
            12'b001010110100: out = 32'b00000000000000111100011000011001;
            12'b001010110101: out = 32'b00000000000000111100010111101110;
            12'b001010110110: out = 32'b00000000000000111100010111000100;
            12'b001010110111: out = 32'b00000000000000111100010110011001;
            12'b001010111000: out = 32'b00000000000000111100010101101111;
            12'b001010111001: out = 32'b00000000000000111100010101000100;
            12'b001010111010: out = 32'b00000000000000111100010100011001;
            12'b001010111011: out = 32'b00000000000000111100010011101110;
            12'b001010111100: out = 32'b00000000000000111100010011000011;
            12'b001010111101: out = 32'b00000000000000111100010010011001;
            12'b001010111110: out = 32'b00000000000000111100010001101110;
            12'b001010111111: out = 32'b00000000000000111100010001000011;
            12'b001011000000: out = 32'b00000000000000111100010000010111;
            12'b001011000001: out = 32'b00000000000000111100001111101100;
            12'b001011000010: out = 32'b00000000000000111100001111000001;
            12'b001011000011: out = 32'b00000000000000111100001110010110;
            12'b001011000100: out = 32'b00000000000000111100001101101010;
            12'b001011000101: out = 32'b00000000000000111100001100111111;
            12'b001011000110: out = 32'b00000000000000111100001100010100;
            12'b001011000111: out = 32'b00000000000000111100001011101000;
            12'b001011001000: out = 32'b00000000000000111100001010111100;
            12'b001011001001: out = 32'b00000000000000111100001010010001;
            12'b001011001010: out = 32'b00000000000000111100001001100101;
            12'b001011001011: out = 32'b00000000000000111100001000111001;
            12'b001011001100: out = 32'b00000000000000111100001000001110;
            12'b001011001101: out = 32'b00000000000000111100000111100010;
            12'b001011001110: out = 32'b00000000000000111100000110110110;
            12'b001011001111: out = 32'b00000000000000111100000110001010;
            12'b001011010000: out = 32'b00000000000000111100000101011110;
            12'b001011010001: out = 32'b00000000000000111100000100110010;
            12'b001011010010: out = 32'b00000000000000111100000100000101;
            12'b001011010011: out = 32'b00000000000000111100000011011001;
            12'b001011010100: out = 32'b00000000000000111100000010101101;
            12'b001011010101: out = 32'b00000000000000111100000010000001;
            12'b001011010110: out = 32'b00000000000000111100000001010100;
            12'b001011010111: out = 32'b00000000000000111100000000101000;
            12'b001011011000: out = 32'b00000000000000111011111111111011;
            12'b001011011001: out = 32'b00000000000000111011111111001111;
            12'b001011011010: out = 32'b00000000000000111011111110100010;
            12'b001011011011: out = 32'b00000000000000111011111101110101;
            12'b001011011100: out = 32'b00000000000000111011111101001001;
            12'b001011011101: out = 32'b00000000000000111011111100011100;
            12'b001011011110: out = 32'b00000000000000111011111011101111;
            12'b001011011111: out = 32'b00000000000000111011111011000010;
            12'b001011100000: out = 32'b00000000000000111011111010010101;
            12'b001011100001: out = 32'b00000000000000111011111001101000;
            12'b001011100010: out = 32'b00000000000000111011111000111011;
            12'b001011100011: out = 32'b00000000000000111011111000001110;
            12'b001011100100: out = 32'b00000000000000111011110111100000;
            12'b001011100101: out = 32'b00000000000000111011110110110011;
            12'b001011100110: out = 32'b00000000000000111011110110000110;
            12'b001011100111: out = 32'b00000000000000111011110101011000;
            12'b001011101000: out = 32'b00000000000000111011110100101011;
            12'b001011101001: out = 32'b00000000000000111011110011111101;
            12'b001011101010: out = 32'b00000000000000111011110011010000;
            12'b001011101011: out = 32'b00000000000000111011110010100010;
            12'b001011101100: out = 32'b00000000000000111011110001110101;
            12'b001011101101: out = 32'b00000000000000111011110001000111;
            12'b001011101110: out = 32'b00000000000000111011110000011001;
            12'b001011101111: out = 32'b00000000000000111011101111101011;
            12'b001011110000: out = 32'b00000000000000111011101110111101;
            12'b001011110001: out = 32'b00000000000000111011101110001111;
            12'b001011110010: out = 32'b00000000000000111011101101100001;
            12'b001011110011: out = 32'b00000000000000111011101100110011;
            12'b001011110100: out = 32'b00000000000000111011101100000101;
            12'b001011110101: out = 32'b00000000000000111011101011010111;
            12'b001011110110: out = 32'b00000000000000111011101010101000;
            12'b001011110111: out = 32'b00000000000000111011101001111010;
            12'b001011111000: out = 32'b00000000000000111011101001001100;
            12'b001011111001: out = 32'b00000000000000111011101000011101;
            12'b001011111010: out = 32'b00000000000000111011100111101111;
            12'b001011111011: out = 32'b00000000000000111011100111000000;
            12'b001011111100: out = 32'b00000000000000111011100110010010;
            12'b001011111101: out = 32'b00000000000000111011100101100011;
            12'b001011111110: out = 32'b00000000000000111011100100110100;
            12'b001011111111: out = 32'b00000000000000111011100100000101;
            12'b001100000000: out = 32'b00000000000000111011100011010110;
            12'b001100000001: out = 32'b00000000000000111011100010101000;
            12'b001100000010: out = 32'b00000000000000111011100001111001;
            12'b001100000011: out = 32'b00000000000000111011100001001010;
            12'b001100000100: out = 32'b00000000000000111011100000011010;
            12'b001100000101: out = 32'b00000000000000111011011111101011;
            12'b001100000110: out = 32'b00000000000000111011011110111100;
            12'b001100000111: out = 32'b00000000000000111011011110001101;
            12'b001100001000: out = 32'b00000000000000111011011101011110;
            12'b001100001001: out = 32'b00000000000000111011011100101110;
            12'b001100001010: out = 32'b00000000000000111011011011111111;
            12'b001100001011: out = 32'b00000000000000111011011011001111;
            12'b001100001100: out = 32'b00000000000000111011011010100000;
            12'b001100001101: out = 32'b00000000000000111011011001110000;
            12'b001100001110: out = 32'b00000000000000111011011001000000;
            12'b001100001111: out = 32'b00000000000000111011011000010001;
            12'b001100010000: out = 32'b00000000000000111011010111100001;
            12'b001100010001: out = 32'b00000000000000111011010110110001;
            12'b001100010010: out = 32'b00000000000000111011010110000001;
            12'b001100010011: out = 32'b00000000000000111011010101010001;
            12'b001100010100: out = 32'b00000000000000111011010100100001;
            12'b001100010101: out = 32'b00000000000000111011010011110001;
            12'b001100010110: out = 32'b00000000000000111011010011000001;
            12'b001100010111: out = 32'b00000000000000111011010010010001;
            12'b001100011000: out = 32'b00000000000000111011010001100001;
            12'b001100011001: out = 32'b00000000000000111011010000110000;
            12'b001100011010: out = 32'b00000000000000111011010000000000;
            12'b001100011011: out = 32'b00000000000000111011001111001111;
            12'b001100011100: out = 32'b00000000000000111011001110011111;
            12'b001100011101: out = 32'b00000000000000111011001101101110;
            12'b001100011110: out = 32'b00000000000000111011001100111110;
            12'b001100011111: out = 32'b00000000000000111011001100001101;
            12'b001100100000: out = 32'b00000000000000111011001011011101;
            12'b001100100001: out = 32'b00000000000000111011001010101100;
            12'b001100100010: out = 32'b00000000000000111011001001111011;
            12'b001100100011: out = 32'b00000000000000111011001001001010;
            12'b001100100100: out = 32'b00000000000000111011001000011001;
            12'b001100100101: out = 32'b00000000000000111011000111101000;
            12'b001100100110: out = 32'b00000000000000111011000110110111;
            12'b001100100111: out = 32'b00000000000000111011000110000110;
            12'b001100101000: out = 32'b00000000000000111011000101010101;
            12'b001100101001: out = 32'b00000000000000111011000100100100;
            12'b001100101010: out = 32'b00000000000000111011000011110010;
            12'b001100101011: out = 32'b00000000000000111011000011000001;
            12'b001100101100: out = 32'b00000000000000111011000010010000;
            12'b001100101101: out = 32'b00000000000000111011000001011110;
            12'b001100101110: out = 32'b00000000000000111011000000101101;
            12'b001100101111: out = 32'b00000000000000111010111111111011;
            12'b001100110000: out = 32'b00000000000000111010111111001001;
            12'b001100110001: out = 32'b00000000000000111010111110011000;
            12'b001100110010: out = 32'b00000000000000111010111101100110;
            12'b001100110011: out = 32'b00000000000000111010111100110100;
            12'b001100110100: out = 32'b00000000000000111010111100000010;
            12'b001100110101: out = 32'b00000000000000111010111011010000;
            12'b001100110110: out = 32'b00000000000000111010111010011110;
            12'b001100110111: out = 32'b00000000000000111010111001101100;
            12'b001100111000: out = 32'b00000000000000111010111000111010;
            12'b001100111001: out = 32'b00000000000000111010111000001000;
            12'b001100111010: out = 32'b00000000000000111010110111010110;
            12'b001100111011: out = 32'b00000000000000111010110110100100;
            12'b001100111100: out = 32'b00000000000000111010110101110001;
            12'b001100111101: out = 32'b00000000000000111010110100111111;
            12'b001100111110: out = 32'b00000000000000111010110100001100;
            12'b001100111111: out = 32'b00000000000000111010110011011010;
            12'b001101000000: out = 32'b00000000000000111010110010100111;
            12'b001101000001: out = 32'b00000000000000111010110001110101;
            12'b001101000010: out = 32'b00000000000000111010110001000010;
            12'b001101000011: out = 32'b00000000000000111010110000001111;
            12'b001101000100: out = 32'b00000000000000111010101111011101;
            12'b001101000101: out = 32'b00000000000000111010101110101010;
            12'b001101000110: out = 32'b00000000000000111010101101110111;
            12'b001101000111: out = 32'b00000000000000111010101101000100;
            12'b001101001000: out = 32'b00000000000000111010101100010001;
            12'b001101001001: out = 32'b00000000000000111010101011011110;
            12'b001101001010: out = 32'b00000000000000111010101010101011;
            12'b001101001011: out = 32'b00000000000000111010101001111000;
            12'b001101001100: out = 32'b00000000000000111010101001000100;
            12'b001101001101: out = 32'b00000000000000111010101000010001;
            12'b001101001110: out = 32'b00000000000000111010100111011110;
            12'b001101001111: out = 32'b00000000000000111010100110101010;
            12'b001101010000: out = 32'b00000000000000111010100101110111;
            12'b001101010001: out = 32'b00000000000000111010100101000011;
            12'b001101010010: out = 32'b00000000000000111010100100010000;
            12'b001101010011: out = 32'b00000000000000111010100011011100;
            12'b001101010100: out = 32'b00000000000000111010100010101000;
            12'b001101010101: out = 32'b00000000000000111010100001110101;
            12'b001101010110: out = 32'b00000000000000111010100001000001;
            12'b001101010111: out = 32'b00000000000000111010100000001101;
            12'b001101011000: out = 32'b00000000000000111010011111011001;
            12'b001101011001: out = 32'b00000000000000111010011110100101;
            12'b001101011010: out = 32'b00000000000000111010011101110001;
            12'b001101011011: out = 32'b00000000000000111010011100111101;
            12'b001101011100: out = 32'b00000000000000111010011100001001;
            12'b001101011101: out = 32'b00000000000000111010011011010100;
            12'b001101011110: out = 32'b00000000000000111010011010100000;
            12'b001101011111: out = 32'b00000000000000111010011001101100;
            12'b001101100000: out = 32'b00000000000000111010011000110111;
            12'b001101100001: out = 32'b00000000000000111010011000000011;
            12'b001101100010: out = 32'b00000000000000111010010111001111;
            12'b001101100011: out = 32'b00000000000000111010010110011010;
            12'b001101100100: out = 32'b00000000000000111010010101100101;
            12'b001101100101: out = 32'b00000000000000111010010100110001;
            12'b001101100110: out = 32'b00000000000000111010010011111100;
            12'b001101100111: out = 32'b00000000000000111010010011000111;
            12'b001101101000: out = 32'b00000000000000111010010010010010;
            12'b001101101001: out = 32'b00000000000000111010010001011101;
            12'b001101101010: out = 32'b00000000000000111010010000101000;
            12'b001101101011: out = 32'b00000000000000111010001111110011;
            12'b001101101100: out = 32'b00000000000000111010001110111110;
            12'b001101101101: out = 32'b00000000000000111010001110001001;
            12'b001101101110: out = 32'b00000000000000111010001101010100;
            12'b001101101111: out = 32'b00000000000000111010001100011111;
            12'b001101110000: out = 32'b00000000000000111010001011101010;
            12'b001101110001: out = 32'b00000000000000111010001010110100;
            12'b001101110010: out = 32'b00000000000000111010001001111111;
            12'b001101110011: out = 32'b00000000000000111010001001001001;
            12'b001101110100: out = 32'b00000000000000111010001000010100;
            12'b001101110101: out = 32'b00000000000000111010000111011110;
            12'b001101110110: out = 32'b00000000000000111010000110101001;
            12'b001101110111: out = 32'b00000000000000111010000101110011;
            12'b001101111000: out = 32'b00000000000000111010000100111101;
            12'b001101111001: out = 32'b00000000000000111010000100000111;
            12'b001101111010: out = 32'b00000000000000111010000011010001;
            12'b001101111011: out = 32'b00000000000000111010000010011100;
            12'b001101111100: out = 32'b00000000000000111010000001100110;
            12'b001101111101: out = 32'b00000000000000111010000000110000;
            12'b001101111110: out = 32'b00000000000000111001111111111001;
            12'b001101111111: out = 32'b00000000000000111001111111000011;
            12'b001110000000: out = 32'b00000000000000111001111110001101;
            12'b001110000001: out = 32'b00000000000000111001111101010111;
            12'b001110000010: out = 32'b00000000000000111001111100100001;
            12'b001110000011: out = 32'b00000000000000111001111011101010;
            12'b001110000100: out = 32'b00000000000000111001111010110100;
            12'b001110000101: out = 32'b00000000000000111001111001111101;
            12'b001110000110: out = 32'b00000000000000111001111001000111;
            12'b001110000111: out = 32'b00000000000000111001111000010000;
            12'b001110001000: out = 32'b00000000000000111001110111011001;
            12'b001110001001: out = 32'b00000000000000111001110110100011;
            12'b001110001010: out = 32'b00000000000000111001110101101100;
            12'b001110001011: out = 32'b00000000000000111001110100110101;
            12'b001110001100: out = 32'b00000000000000111001110011111110;
            12'b001110001101: out = 32'b00000000000000111001110011000111;
            12'b001110001110: out = 32'b00000000000000111001110010010000;
            12'b001110001111: out = 32'b00000000000000111001110001011001;
            12'b001110010000: out = 32'b00000000000000111001110000100010;
            12'b001110010001: out = 32'b00000000000000111001101111101011;
            12'b001110010010: out = 32'b00000000000000111001101110110100;
            12'b001110010011: out = 32'b00000000000000111001101101111101;
            12'b001110010100: out = 32'b00000000000000111001101101000101;
            12'b001110010101: out = 32'b00000000000000111001101100001110;
            12'b001110010110: out = 32'b00000000000000111001101011010110;
            12'b001110010111: out = 32'b00000000000000111001101010011111;
            12'b001110011000: out = 32'b00000000000000111001101001100111;
            12'b001110011001: out = 32'b00000000000000111001101000110000;
            12'b001110011010: out = 32'b00000000000000111001100111111000;
            12'b001110011011: out = 32'b00000000000000111001100111000000;
            12'b001110011100: out = 32'b00000000000000111001100110001001;
            12'b001110011101: out = 32'b00000000000000111001100101010001;
            12'b001110011110: out = 32'b00000000000000111001100100011001;
            12'b001110011111: out = 32'b00000000000000111001100011100001;
            12'b001110100000: out = 32'b00000000000000111001100010101001;
            12'b001110100001: out = 32'b00000000000000111001100001110001;
            12'b001110100010: out = 32'b00000000000000111001100000111001;
            12'b001110100011: out = 32'b00000000000000111001100000000000;
            12'b001110100100: out = 32'b00000000000000111001011111001000;
            12'b001110100101: out = 32'b00000000000000111001011110010000;
            12'b001110100110: out = 32'b00000000000000111001011101011000;
            12'b001110100111: out = 32'b00000000000000111001011100011111;
            12'b001110101000: out = 32'b00000000000000111001011011100111;
            12'b001110101001: out = 32'b00000000000000111001011010101110;
            12'b001110101010: out = 32'b00000000000000111001011001110110;
            12'b001110101011: out = 32'b00000000000000111001011000111101;
            12'b001110101100: out = 32'b00000000000000111001011000000100;
            12'b001110101101: out = 32'b00000000000000111001010111001100;
            12'b001110101110: out = 32'b00000000000000111001010110010011;
            12'b001110101111: out = 32'b00000000000000111001010101011010;
            12'b001110110000: out = 32'b00000000000000111001010100100001;
            12'b001110110001: out = 32'b00000000000000111001010011101000;
            12'b001110110010: out = 32'b00000000000000111001010010101111;
            12'b001110110011: out = 32'b00000000000000111001010001110110;
            12'b001110110100: out = 32'b00000000000000111001010000111101;
            12'b001110110101: out = 32'b00000000000000111001010000000100;
            12'b001110110110: out = 32'b00000000000000111001001111001010;
            12'b001110110111: out = 32'b00000000000000111001001110010001;
            12'b001110111000: out = 32'b00000000000000111001001101011000;
            12'b001110111001: out = 32'b00000000000000111001001100011110;
            12'b001110111010: out = 32'b00000000000000111001001011100101;
            12'b001110111011: out = 32'b00000000000000111001001010101011;
            12'b001110111100: out = 32'b00000000000000111001001001110010;
            12'b001110111101: out = 32'b00000000000000111001001000111000;
            12'b001110111110: out = 32'b00000000000000111001000111111111;
            12'b001110111111: out = 32'b00000000000000111001000111000101;
            12'b001111000000: out = 32'b00000000000000111001000110001011;
            12'b001111000001: out = 32'b00000000000000111001000101010001;
            12'b001111000010: out = 32'b00000000000000111001000100010111;
            12'b001111000011: out = 32'b00000000000000111001000011011101;
            12'b001111000100: out = 32'b00000000000000111001000010100011;
            12'b001111000101: out = 32'b00000000000000111001000001101001;
            12'b001111000110: out = 32'b00000000000000111001000000101111;
            12'b001111000111: out = 32'b00000000000000111000111111110101;
            12'b001111001000: out = 32'b00000000000000111000111110111011;
            12'b001111001001: out = 32'b00000000000000111000111110000000;
            12'b001111001010: out = 32'b00000000000000111000111101000110;
            12'b001111001011: out = 32'b00000000000000111000111100001100;
            12'b001111001100: out = 32'b00000000000000111000111011010001;
            12'b001111001101: out = 32'b00000000000000111000111010010111;
            12'b001111001110: out = 32'b00000000000000111000111001011100;
            12'b001111001111: out = 32'b00000000000000111000111000100001;
            12'b001111010000: out = 32'b00000000000000111000110111100111;
            12'b001111010001: out = 32'b00000000000000111000110110101100;
            12'b001111010010: out = 32'b00000000000000111000110101110001;
            12'b001111010011: out = 32'b00000000000000111000110100110110;
            12'b001111010100: out = 32'b00000000000000111000110011111011;
            12'b001111010101: out = 32'b00000000000000111000110011000000;
            12'b001111010110: out = 32'b00000000000000111000110010000101;
            12'b001111010111: out = 32'b00000000000000111000110001001010;
            12'b001111011000: out = 32'b00000000000000111000110000001111;
            12'b001111011001: out = 32'b00000000000000111000101111010100;
            12'b001111011010: out = 32'b00000000000000111000101110011001;
            12'b001111011011: out = 32'b00000000000000111000101101011101;
            12'b001111011100: out = 32'b00000000000000111000101100100010;
            12'b001111011101: out = 32'b00000000000000111000101011100111;
            12'b001111011110: out = 32'b00000000000000111000101010101011;
            12'b001111011111: out = 32'b00000000000000111000101001110000;
            12'b001111100000: out = 32'b00000000000000111000101000110100;
            12'b001111100001: out = 32'b00000000000000111000100111111000;
            12'b001111100010: out = 32'b00000000000000111000100110111101;
            12'b001111100011: out = 32'b00000000000000111000100110000001;
            12'b001111100100: out = 32'b00000000000000111000100101000101;
            12'b001111100101: out = 32'b00000000000000111000100100001001;
            12'b001111100110: out = 32'b00000000000000111000100011001101;
            12'b001111100111: out = 32'b00000000000000111000100010010001;
            12'b001111101000: out = 32'b00000000000000111000100001010101;
            12'b001111101001: out = 32'b00000000000000111000100000011001;
            12'b001111101010: out = 32'b00000000000000111000011111011101;
            12'b001111101011: out = 32'b00000000000000111000011110100001;
            12'b001111101100: out = 32'b00000000000000111000011101100101;
            12'b001111101101: out = 32'b00000000000000111000011100101001;
            12'b001111101110: out = 32'b00000000000000111000011011101100;
            12'b001111101111: out = 32'b00000000000000111000011010110000;
            12'b001111110000: out = 32'b00000000000000111000011001110011;
            12'b001111110001: out = 32'b00000000000000111000011000110111;
            12'b001111110010: out = 32'b00000000000000111000010111111010;
            12'b001111110011: out = 32'b00000000000000111000010110111110;
            12'b001111110100: out = 32'b00000000000000111000010110000001;
            12'b001111110101: out = 32'b00000000000000111000010101000100;
            12'b001111110110: out = 32'b00000000000000111000010100000111;
            12'b001111110111: out = 32'b00000000000000111000010011001011;
            12'b001111111000: out = 32'b00000000000000111000010010001110;
            12'b001111111001: out = 32'b00000000000000111000010001010001;
            12'b001111111010: out = 32'b00000000000000111000010000010100;
            12'b001111111011: out = 32'b00000000000000111000001111010111;
            12'b001111111100: out = 32'b00000000000000111000001110011010;
            12'b001111111101: out = 32'b00000000000000111000001101011100;
            12'b001111111110: out = 32'b00000000000000111000001100011111;
            12'b001111111111: out = 32'b00000000000000111000001011100010;
            12'b010000000000: out = 32'b00000000000000111000001010100101;
            12'b010000000001: out = 32'b00000000000000111000001001100111;
            12'b010000000010: out = 32'b00000000000000111000001000101010;
            12'b010000000011: out = 32'b00000000000000111000000111101100;
            12'b010000000100: out = 32'b00000000000000111000000110101111;
            12'b010000000101: out = 32'b00000000000000111000000101110001;
            12'b010000000110: out = 32'b00000000000000111000000100110011;
            12'b010000000111: out = 32'b00000000000000111000000011110110;
            12'b010000001000: out = 32'b00000000000000111000000010111000;
            12'b010000001001: out = 32'b00000000000000111000000001111010;
            12'b010000001010: out = 32'b00000000000000111000000000111100;
            12'b010000001011: out = 32'b00000000000000110111111111111110;
            12'b010000001100: out = 32'b00000000000000110111111111000000;
            12'b010000001101: out = 32'b00000000000000110111111110000010;
            12'b010000001110: out = 32'b00000000000000110111111101000100;
            12'b010000001111: out = 32'b00000000000000110111111100000110;
            12'b010000010000: out = 32'b00000000000000110111111011001000;
            12'b010000010001: out = 32'b00000000000000110111111010001001;
            12'b010000010010: out = 32'b00000000000000110111111001001011;
            12'b010000010011: out = 32'b00000000000000110111111000001101;
            12'b010000010100: out = 32'b00000000000000110111110111001110;
            12'b010000010101: out = 32'b00000000000000110111110110010000;
            12'b010000010110: out = 32'b00000000000000110111110101010001;
            12'b010000010111: out = 32'b00000000000000110111110100010011;
            12'b010000011000: out = 32'b00000000000000110111110011010100;
            12'b010000011001: out = 32'b00000000000000110111110010010101;
            12'b010000011010: out = 32'b00000000000000110111110001010110;
            12'b010000011011: out = 32'b00000000000000110111110000011000;
            12'b010000011100: out = 32'b00000000000000110111101111011001;
            12'b010000011101: out = 32'b00000000000000110111101110011010;
            12'b010000011110: out = 32'b00000000000000110111101101011011;
            12'b010000011111: out = 32'b00000000000000110111101100011100;
            12'b010000100000: out = 32'b00000000000000110111101011011101;
            12'b010000100001: out = 32'b00000000000000110111101010011110;
            12'b010000100010: out = 32'b00000000000000110111101001011110;
            12'b010000100011: out = 32'b00000000000000110111101000011111;
            12'b010000100100: out = 32'b00000000000000110111100111100000;
            12'b010000100101: out = 32'b00000000000000110111100110100001;
            12'b010000100110: out = 32'b00000000000000110111100101100001;
            12'b010000100111: out = 32'b00000000000000110111100100100010;
            12'b010000101000: out = 32'b00000000000000110111100011100010;
            12'b010000101001: out = 32'b00000000000000110111100010100011;
            12'b010000101010: out = 32'b00000000000000110111100001100011;
            12'b010000101011: out = 32'b00000000000000110111100000100011;
            12'b010000101100: out = 32'b00000000000000110111011111100011;
            12'b010000101101: out = 32'b00000000000000110111011110100100;
            12'b010000101110: out = 32'b00000000000000110111011101100100;
            12'b010000101111: out = 32'b00000000000000110111011100100100;
            12'b010000110000: out = 32'b00000000000000110111011011100100;
            12'b010000110001: out = 32'b00000000000000110111011010100100;
            12'b010000110010: out = 32'b00000000000000110111011001100100;
            12'b010000110011: out = 32'b00000000000000110111011000100100;
            12'b010000110100: out = 32'b00000000000000110111010111100100;
            12'b010000110101: out = 32'b00000000000000110111010110100011;
            12'b010000110110: out = 32'b00000000000000110111010101100011;
            12'b010000110111: out = 32'b00000000000000110111010100100011;
            12'b010000111000: out = 32'b00000000000000110111010011100010;
            12'b010000111001: out = 32'b00000000000000110111010010100010;
            12'b010000111010: out = 32'b00000000000000110111010001100001;
            12'b010000111011: out = 32'b00000000000000110111010000100001;
            12'b010000111100: out = 32'b00000000000000110111001111100000;
            12'b010000111101: out = 32'b00000000000000110111001110100000;
            12'b010000111110: out = 32'b00000000000000110111001101011111;
            12'b010000111111: out = 32'b00000000000000110111001100011110;
            12'b010001000000: out = 32'b00000000000000110111001011011101;
            12'b010001000001: out = 32'b00000000000000110111001010011100;
            12'b010001000010: out = 32'b00000000000000110111001001011100;
            12'b010001000011: out = 32'b00000000000000110111001000011011;
            12'b010001000100: out = 32'b00000000000000110111000111011010;
            12'b010001000101: out = 32'b00000000000000110111000110011000;
            12'b010001000110: out = 32'b00000000000000110111000101010111;
            12'b010001000111: out = 32'b00000000000000110111000100010110;
            12'b010001001000: out = 32'b00000000000000110111000011010101;
            12'b010001001001: out = 32'b00000000000000110111000010010100;
            12'b010001001010: out = 32'b00000000000000110111000001010010;
            12'b010001001011: out = 32'b00000000000000110111000000010001;
            12'b010001001100: out = 32'b00000000000000110110111111001111;
            12'b010001001101: out = 32'b00000000000000110110111110001110;
            12'b010001001110: out = 32'b00000000000000110110111101001100;
            12'b010001001111: out = 32'b00000000000000110110111100001011;
            12'b010001010000: out = 32'b00000000000000110110111011001001;
            12'b010001010001: out = 32'b00000000000000110110111010000111;
            12'b010001010010: out = 32'b00000000000000110110111001000101;
            12'b010001010011: out = 32'b00000000000000110110111000000100;
            12'b010001010100: out = 32'b00000000000000110110110111000010;
            12'b010001010101: out = 32'b00000000000000110110110110000000;
            12'b010001010110: out = 32'b00000000000000110110110100111110;
            12'b010001010111: out = 32'b00000000000000110110110011111100;
            12'b010001011000: out = 32'b00000000000000110110110010111010;
            12'b010001011001: out = 32'b00000000000000110110110001110111;
            12'b010001011010: out = 32'b00000000000000110110110000110101;
            12'b010001011011: out = 32'b00000000000000110110101111110011;
            12'b010001011100: out = 32'b00000000000000110110101110110001;
            12'b010001011101: out = 32'b00000000000000110110101101101110;
            12'b010001011110: out = 32'b00000000000000110110101100101100;
            12'b010001011111: out = 32'b00000000000000110110101011101001;
            12'b010001100000: out = 32'b00000000000000110110101010100111;
            12'b010001100001: out = 32'b00000000000000110110101001100100;
            12'b010001100010: out = 32'b00000000000000110110101000100010;
            12'b010001100011: out = 32'b00000000000000110110100111011111;
            12'b010001100100: out = 32'b00000000000000110110100110011100;
            12'b010001100101: out = 32'b00000000000000110110100101011001;
            12'b010001100110: out = 32'b00000000000000110110100100010110;
            12'b010001100111: out = 32'b00000000000000110110100011010100;
            12'b010001101000: out = 32'b00000000000000110110100010010001;
            12'b010001101001: out = 32'b00000000000000110110100001001110;
            12'b010001101010: out = 32'b00000000000000110110100000001010;
            12'b010001101011: out = 32'b00000000000000110110011111000111;
            12'b010001101100: out = 32'b00000000000000110110011110000100;
            12'b010001101101: out = 32'b00000000000000110110011101000001;
            12'b010001101110: out = 32'b00000000000000110110011011111110;
            12'b010001101111: out = 32'b00000000000000110110011010111010;
            12'b010001110000: out = 32'b00000000000000110110011001110111;
            12'b010001110001: out = 32'b00000000000000110110011000110100;
            12'b010001110010: out = 32'b00000000000000110110010111110000;
            12'b010001110011: out = 32'b00000000000000110110010110101100;
            12'b010001110100: out = 32'b00000000000000110110010101101001;
            12'b010001110101: out = 32'b00000000000000110110010100100101;
            12'b010001110110: out = 32'b00000000000000110110010011100010;
            12'b010001110111: out = 32'b00000000000000110110010010011110;
            12'b010001111000: out = 32'b00000000000000110110010001011010;
            12'b010001111001: out = 32'b00000000000000110110010000010110;
            12'b010001111010: out = 32'b00000000000000110110001111010010;
            12'b010001111011: out = 32'b00000000000000110110001110001110;
            12'b010001111100: out = 32'b00000000000000110110001101001010;
            12'b010001111101: out = 32'b00000000000000110110001100000110;
            12'b010001111110: out = 32'b00000000000000110110001011000010;
            12'b010001111111: out = 32'b00000000000000110110001001111110;
            12'b010010000000: out = 32'b00000000000000110110001000111010;
            12'b010010000001: out = 32'b00000000000000110110000111110101;
            12'b010010000010: out = 32'b00000000000000110110000110110001;
            12'b010010000011: out = 32'b00000000000000110110000101101101;
            12'b010010000100: out = 32'b00000000000000110110000100101000;
            12'b010010000101: out = 32'b00000000000000110110000011100100;
            12'b010010000110: out = 32'b00000000000000110110000010011111;
            12'b010010000111: out = 32'b00000000000000110110000001011010;
            12'b010010001000: out = 32'b00000000000000110110000000010110;
            12'b010010001001: out = 32'b00000000000000110101111111010001;
            12'b010010001010: out = 32'b00000000000000110101111110001100;
            12'b010010001011: out = 32'b00000000000000110101111101000111;
            12'b010010001100: out = 32'b00000000000000110101111100000011;
            12'b010010001101: out = 32'b00000000000000110101111010111110;
            12'b010010001110: out = 32'b00000000000000110101111001111001;
            12'b010010001111: out = 32'b00000000000000110101111000110100;
            12'b010010010000: out = 32'b00000000000000110101110111101111;
            12'b010010010001: out = 32'b00000000000000110101110110101001;
            12'b010010010010: out = 32'b00000000000000110101110101100100;
            12'b010010010011: out = 32'b00000000000000110101110100011111;
            12'b010010010100: out = 32'b00000000000000110101110011011010;
            12'b010010010101: out = 32'b00000000000000110101110010010100;
            12'b010010010110: out = 32'b00000000000000110101110001001111;
            12'b010010010111: out = 32'b00000000000000110101110000001010;
            12'b010010011000: out = 32'b00000000000000110101101111000100;
            12'b010010011001: out = 32'b00000000000000110101101101111110;
            12'b010010011010: out = 32'b00000000000000110101101100111001;
            12'b010010011011: out = 32'b00000000000000110101101011110011;
            12'b010010011100: out = 32'b00000000000000110101101010101110;
            12'b010010011101: out = 32'b00000000000000110101101001101000;
            12'b010010011110: out = 32'b00000000000000110101101000100010;
            12'b010010011111: out = 32'b00000000000000110101100111011100;
            12'b010010100000: out = 32'b00000000000000110101100110010110;
            12'b010010100001: out = 32'b00000000000000110101100101010000;
            12'b010010100010: out = 32'b00000000000000110101100100001010;
            12'b010010100011: out = 32'b00000000000000110101100011000100;
            12'b010010100100: out = 32'b00000000000000110101100001111110;
            12'b010010100101: out = 32'b00000000000000110101100000111000;
            12'b010010100110: out = 32'b00000000000000110101011111110010;
            12'b010010100111: out = 32'b00000000000000110101011110101011;
            12'b010010101000: out = 32'b00000000000000110101011101100101;
            12'b010010101001: out = 32'b00000000000000110101011100011111;
            12'b010010101010: out = 32'b00000000000000110101011011011000;
            12'b010010101011: out = 32'b00000000000000110101011010010010;
            12'b010010101100: out = 32'b00000000000000110101011001001011;
            12'b010010101101: out = 32'b00000000000000110101011000000100;
            12'b010010101110: out = 32'b00000000000000110101010110111110;
            12'b010010101111: out = 32'b00000000000000110101010101110111;
            12'b010010110000: out = 32'b00000000000000110101010100110000;
            12'b010010110001: out = 32'b00000000000000110101010011101010;
            12'b010010110010: out = 32'b00000000000000110101010010100011;
            12'b010010110011: out = 32'b00000000000000110101010001011100;
            12'b010010110100: out = 32'b00000000000000110101010000010101;
            12'b010010110101: out = 32'b00000000000000110101001111001110;
            12'b010010110110: out = 32'b00000000000000110101001110000111;
            12'b010010110111: out = 32'b00000000000000110101001101000000;
            12'b010010111000: out = 32'b00000000000000110101001011111000;
            12'b010010111001: out = 32'b00000000000000110101001010110001;
            12'b010010111010: out = 32'b00000000000000110101001001101010;
            12'b010010111011: out = 32'b00000000000000110101001000100011;
            12'b010010111100: out = 32'b00000000000000110101000111011011;
            12'b010010111101: out = 32'b00000000000000110101000110010100;
            12'b010010111110: out = 32'b00000000000000110101000101001100;
            12'b010010111111: out = 32'b00000000000000110101000100000101;
            12'b010011000000: out = 32'b00000000000000110101000010111101;
            12'b010011000001: out = 32'b00000000000000110101000001110110;
            12'b010011000010: out = 32'b00000000000000110101000000101110;
            12'b010011000011: out = 32'b00000000000000110100111111100110;
            12'b010011000100: out = 32'b00000000000000110100111110011110;
            12'b010011000101: out = 32'b00000000000000110100111101010110;
            12'b010011000110: out = 32'b00000000000000110100111100001111;
            12'b010011000111: out = 32'b00000000000000110100111011000111;
            12'b010011001000: out = 32'b00000000000000110100111001111111;
            12'b010011001001: out = 32'b00000000000000110100111000110111;
            12'b010011001010: out = 32'b00000000000000110100110111101110;
            12'b010011001011: out = 32'b00000000000000110100110110100110;
            12'b010011001100: out = 32'b00000000000000110100110101011110;
            12'b010011001101: out = 32'b00000000000000110100110100010110;
            12'b010011001110: out = 32'b00000000000000110100110011001110;
            12'b010011001111: out = 32'b00000000000000110100110010000101;
            12'b010011010000: out = 32'b00000000000000110100110000111101;
            12'b010011010001: out = 32'b00000000000000110100101111110100;
            12'b010011010010: out = 32'b00000000000000110100101110101100;
            12'b010011010011: out = 32'b00000000000000110100101101100011;
            12'b010011010100: out = 32'b00000000000000110100101100011011;
            12'b010011010101: out = 32'b00000000000000110100101011010010;
            12'b010011010110: out = 32'b00000000000000110100101010001001;
            12'b010011010111: out = 32'b00000000000000110100101001000000;
            12'b010011011000: out = 32'b00000000000000110100100111111000;
            12'b010011011001: out = 32'b00000000000000110100100110101111;
            12'b010011011010: out = 32'b00000000000000110100100101100110;
            12'b010011011011: out = 32'b00000000000000110100100100011101;
            12'b010011011100: out = 32'b00000000000000110100100011010100;
            12'b010011011101: out = 32'b00000000000000110100100010001011;
            12'b010011011110: out = 32'b00000000000000110100100001000010;
            12'b010011011111: out = 32'b00000000000000110100011111111000;
            12'b010011100000: out = 32'b00000000000000110100011110101111;
            12'b010011100001: out = 32'b00000000000000110100011101100110;
            12'b010011100010: out = 32'b00000000000000110100011100011101;
            12'b010011100011: out = 32'b00000000000000110100011011010011;
            12'b010011100100: out = 32'b00000000000000110100011010001010;
            12'b010011100101: out = 32'b00000000000000110100011001000000;
            12'b010011100110: out = 32'b00000000000000110100010111110111;
            12'b010011100111: out = 32'b00000000000000110100010110101101;
            12'b010011101000: out = 32'b00000000000000110100010101100011;
            12'b010011101001: out = 32'b00000000000000110100010100011010;
            12'b010011101010: out = 32'b00000000000000110100010011010000;
            12'b010011101011: out = 32'b00000000000000110100010010000110;
            12'b010011101100: out = 32'b00000000000000110100010000111100;
            12'b010011101101: out = 32'b00000000000000110100001111110010;
            12'b010011101110: out = 32'b00000000000000110100001110101000;
            12'b010011101111: out = 32'b00000000000000110100001101011110;
            12'b010011110000: out = 32'b00000000000000110100001100010100;
            12'b010011110001: out = 32'b00000000000000110100001011001010;
            12'b010011110010: out = 32'b00000000000000110100001010000000;
            12'b010011110011: out = 32'b00000000000000110100001000110110;
            12'b010011110100: out = 32'b00000000000000110100000111101100;
            12'b010011110101: out = 32'b00000000000000110100000110100001;
            12'b010011110110: out = 32'b00000000000000110100000101010111;
            12'b010011110111: out = 32'b00000000000000110100000100001101;
            12'b010011111000: out = 32'b00000000000000110100000011000010;
            12'b010011111001: out = 32'b00000000000000110100000001111000;
            12'b010011111010: out = 32'b00000000000000110100000000101101;
            12'b010011111011: out = 32'b00000000000000110011111111100010;
            12'b010011111100: out = 32'b00000000000000110011111110011000;
            12'b010011111101: out = 32'b00000000000000110011111101001101;
            12'b010011111110: out = 32'b00000000000000110011111100000010;
            12'b010011111111: out = 32'b00000000000000110011111010110111;
            12'b010100000000: out = 32'b00000000000000110011111001101101;
            12'b010100000001: out = 32'b00000000000000110011111000100010;
            12'b010100000010: out = 32'b00000000000000110011110111010111;
            12'b010100000011: out = 32'b00000000000000110011110110001100;
            12'b010100000100: out = 32'b00000000000000110011110101000001;
            12'b010100000101: out = 32'b00000000000000110011110011110110;
            12'b010100000110: out = 32'b00000000000000110011110010101010;
            12'b010100000111: out = 32'b00000000000000110011110001011111;
            12'b010100001000: out = 32'b00000000000000110011110000010100;
            12'b010100001001: out = 32'b00000000000000110011101111001001;
            12'b010100001010: out = 32'b00000000000000110011101101111101;
            12'b010100001011: out = 32'b00000000000000110011101100110010;
            12'b010100001100: out = 32'b00000000000000110011101011100110;
            12'b010100001101: out = 32'b00000000000000110011101010011011;
            12'b010100001110: out = 32'b00000000000000110011101001001111;
            12'b010100001111: out = 32'b00000000000000110011101000000100;
            12'b010100010000: out = 32'b00000000000000110011100110111000;
            12'b010100010001: out = 32'b00000000000000110011100101101100;
            12'b010100010010: out = 32'b00000000000000110011100100100000;
            12'b010100010011: out = 32'b00000000000000110011100011010101;
            12'b010100010100: out = 32'b00000000000000110011100010001001;
            12'b010100010101: out = 32'b00000000000000110011100000111101;
            12'b010100010110: out = 32'b00000000000000110011011111110001;
            12'b010100010111: out = 32'b00000000000000110011011110100101;
            12'b010100011000: out = 32'b00000000000000110011011101011001;
            12'b010100011001: out = 32'b00000000000000110011011100001101;
            12'b010100011010: out = 32'b00000000000000110011011011000000;
            12'b010100011011: out = 32'b00000000000000110011011001110100;
            12'b010100011100: out = 32'b00000000000000110011011000101000;
            12'b010100011101: out = 32'b00000000000000110011010111011011;
            12'b010100011110: out = 32'b00000000000000110011010110001111;
            12'b010100011111: out = 32'b00000000000000110011010101000011;
            12'b010100100000: out = 32'b00000000000000110011010011110110;
            12'b010100100001: out = 32'b00000000000000110011010010101010;
            12'b010100100010: out = 32'b00000000000000110011010001011101;
            12'b010100100011: out = 32'b00000000000000110011010000010000;
            12'b010100100100: out = 32'b00000000000000110011001111000100;
            12'b010100100101: out = 32'b00000000000000110011001101110111;
            12'b010100100110: out = 32'b00000000000000110011001100101010;
            12'b010100100111: out = 32'b00000000000000110011001011011101;
            12'b010100101000: out = 32'b00000000000000110011001010010001;
            12'b010100101001: out = 32'b00000000000000110011001001000100;
            12'b010100101010: out = 32'b00000000000000110011000111110111;
            12'b010100101011: out = 32'b00000000000000110011000110101010;
            12'b010100101100: out = 32'b00000000000000110011000101011101;
            12'b010100101101: out = 32'b00000000000000110011000100001111;
            12'b010100101110: out = 32'b00000000000000110011000011000010;
            12'b010100101111: out = 32'b00000000000000110011000001110101;
            12'b010100110000: out = 32'b00000000000000110011000000101000;
            12'b010100110001: out = 32'b00000000000000110010111111011010;
            12'b010100110010: out = 32'b00000000000000110010111110001101;
            12'b010100110011: out = 32'b00000000000000110010111101000000;
            12'b010100110100: out = 32'b00000000000000110010111011110010;
            12'b010100110101: out = 32'b00000000000000110010111010100101;
            12'b010100110110: out = 32'b00000000000000110010111001010111;
            12'b010100110111: out = 32'b00000000000000110010111000001001;
            12'b010100111000: out = 32'b00000000000000110010110110111100;
            12'b010100111001: out = 32'b00000000000000110010110101101110;
            12'b010100111010: out = 32'b00000000000000110010110100100000;
            12'b010100111011: out = 32'b00000000000000110010110011010010;
            12'b010100111100: out = 32'b00000000000000110010110010000100;
            12'b010100111101: out = 32'b00000000000000110010110000110111;
            12'b010100111110: out = 32'b00000000000000110010101111101001;
            12'b010100111111: out = 32'b00000000000000110010101110011011;
            12'b010101000000: out = 32'b00000000000000110010101101001100;
            12'b010101000001: out = 32'b00000000000000110010101011111110;
            12'b010101000010: out = 32'b00000000000000110010101010110000;
            12'b010101000011: out = 32'b00000000000000110010101001100010;
            12'b010101000100: out = 32'b00000000000000110010101000010100;
            12'b010101000101: out = 32'b00000000000000110010100111000101;
            12'b010101000110: out = 32'b00000000000000110010100101110111;
            12'b010101000111: out = 32'b00000000000000110010100100101001;
            12'b010101001000: out = 32'b00000000000000110010100011011010;
            12'b010101001001: out = 32'b00000000000000110010100010001100;
            12'b010101001010: out = 32'b00000000000000110010100000111101;
            12'b010101001011: out = 32'b00000000000000110010011111101110;
            12'b010101001100: out = 32'b00000000000000110010011110100000;
            12'b010101001101: out = 32'b00000000000000110010011101010001;
            12'b010101001110: out = 32'b00000000000000110010011100000010;
            12'b010101001111: out = 32'b00000000000000110010011010110011;
            12'b010101010000: out = 32'b00000000000000110010011001100101;
            12'b010101010001: out = 32'b00000000000000110010011000010110;
            12'b010101010010: out = 32'b00000000000000110010010111000111;
            12'b010101010011: out = 32'b00000000000000110010010101111000;
            12'b010101010100: out = 32'b00000000000000110010010100101001;
            12'b010101010101: out = 32'b00000000000000110010010011011010;
            12'b010101010110: out = 32'b00000000000000110010010010001010;
            12'b010101010111: out = 32'b00000000000000110010010000111011;
            12'b010101011000: out = 32'b00000000000000110010001111101100;
            12'b010101011001: out = 32'b00000000000000110010001110011101;
            12'b010101011010: out = 32'b00000000000000110010001101001101;
            12'b010101011011: out = 32'b00000000000000110010001011111110;
            12'b010101011100: out = 32'b00000000000000110010001010101110;
            12'b010101011101: out = 32'b00000000000000110010001001011111;
            12'b010101011110: out = 32'b00000000000000110010001000001111;
            12'b010101011111: out = 32'b00000000000000110010000111000000;
            12'b010101100000: out = 32'b00000000000000110010000101110000;
            12'b010101100001: out = 32'b00000000000000110010000100100000;
            12'b010101100010: out = 32'b00000000000000110010000011010001;
            12'b010101100011: out = 32'b00000000000000110010000010000001;
            12'b010101100100: out = 32'b00000000000000110010000000110001;
            12'b010101100101: out = 32'b00000000000000110001111111100001;
            12'b010101100110: out = 32'b00000000000000110001111110010001;
            12'b010101100111: out = 32'b00000000000000110001111101000001;
            12'b010101101000: out = 32'b00000000000000110001111011110001;
            12'b010101101001: out = 32'b00000000000000110001111010100001;
            12'b010101101010: out = 32'b00000000000000110001111001010001;
            12'b010101101011: out = 32'b00000000000000110001111000000001;
            12'b010101101100: out = 32'b00000000000000110001110110110000;
            12'b010101101101: out = 32'b00000000000000110001110101100000;
            12'b010101101110: out = 32'b00000000000000110001110100010000;
            12'b010101101111: out = 32'b00000000000000110001110010111111;
            12'b010101110000: out = 32'b00000000000000110001110001101111;
            12'b010101110001: out = 32'b00000000000000110001110000011111;
            12'b010101110010: out = 32'b00000000000000110001101111001110;
            12'b010101110011: out = 32'b00000000000000110001101101111101;
            12'b010101110100: out = 32'b00000000000000110001101100101101;
            12'b010101110101: out = 32'b00000000000000110001101011011100;
            12'b010101110110: out = 32'b00000000000000110001101010001011;
            12'b010101110111: out = 32'b00000000000000110001101000111011;
            12'b010101111000: out = 32'b00000000000000110001100111101010;
            12'b010101111001: out = 32'b00000000000000110001100110011001;
            12'b010101111010: out = 32'b00000000000000110001100101001000;
            12'b010101111011: out = 32'b00000000000000110001100011110111;
            12'b010101111100: out = 32'b00000000000000110001100010100110;
            12'b010101111101: out = 32'b00000000000000110001100001010101;
            12'b010101111110: out = 32'b00000000000000110001100000000100;
            12'b010101111111: out = 32'b00000000000000110001011110110011;
            12'b010110000000: out = 32'b00000000000000110001011101100010;
            12'b010110000001: out = 32'b00000000000000110001011100010000;
            12'b010110000010: out = 32'b00000000000000110001011010111111;
            12'b010110000011: out = 32'b00000000000000110001011001101110;
            12'b010110000100: out = 32'b00000000000000110001011000011100;
            12'b010110000101: out = 32'b00000000000000110001010111001011;
            12'b010110000110: out = 32'b00000000000000110001010101111001;
            12'b010110000111: out = 32'b00000000000000110001010100101000;
            12'b010110001000: out = 32'b00000000000000110001010011010110;
            12'b010110001001: out = 32'b00000000000000110001010010000101;
            12'b010110001010: out = 32'b00000000000000110001010000110011;
            12'b010110001011: out = 32'b00000000000000110001001111100001;
            12'b010110001100: out = 32'b00000000000000110001001110001111;
            12'b010110001101: out = 32'b00000000000000110001001100111101;
            12'b010110001110: out = 32'b00000000000000110001001011101100;
            12'b010110001111: out = 32'b00000000000000110001001010011010;
            12'b010110010000: out = 32'b00000000000000110001001001001000;
            12'b010110010001: out = 32'b00000000000000110001000111110110;
            12'b010110010010: out = 32'b00000000000000110001000110100100;
            12'b010110010011: out = 32'b00000000000000110001000101010001;
            12'b010110010100: out = 32'b00000000000000110001000011111111;
            12'b010110010101: out = 32'b00000000000000110001000010101101;
            12'b010110010110: out = 32'b00000000000000110001000001011011;
            12'b010110010111: out = 32'b00000000000000110001000000001001;
            12'b010110011000: out = 32'b00000000000000110000111110110110;
            12'b010110011001: out = 32'b00000000000000110000111101100100;
            12'b010110011010: out = 32'b00000000000000110000111100010001;
            12'b010110011011: out = 32'b00000000000000110000111010111111;
            12'b010110011100: out = 32'b00000000000000110000111001101100;
            12'b010110011101: out = 32'b00000000000000110000111000011010;
            12'b010110011110: out = 32'b00000000000000110000110111000111;
            12'b010110011111: out = 32'b00000000000000110000110101110100;
            12'b010110100000: out = 32'b00000000000000110000110100100010;
            12'b010110100001: out = 32'b00000000000000110000110011001111;
            12'b010110100010: out = 32'b00000000000000110000110001111100;
            12'b010110100011: out = 32'b00000000000000110000110000101001;
            12'b010110100100: out = 32'b00000000000000110000101111010110;
            12'b010110100101: out = 32'b00000000000000110000101110000011;
            12'b010110100110: out = 32'b00000000000000110000101100110000;
            12'b010110100111: out = 32'b00000000000000110000101011011101;
            12'b010110101000: out = 32'b00000000000000110000101010001010;
            12'b010110101001: out = 32'b00000000000000110000101000110111;
            12'b010110101010: out = 32'b00000000000000110000100111100100;
            12'b010110101011: out = 32'b00000000000000110000100110010000;
            12'b010110101100: out = 32'b00000000000000110000100100111101;
            12'b010110101101: out = 32'b00000000000000110000100011101010;
            12'b010110101110: out = 32'b00000000000000110000100010010110;
            12'b010110101111: out = 32'b00000000000000110000100001000011;
            12'b010110110000: out = 32'b00000000000000110000011111101111;
            12'b010110110001: out = 32'b00000000000000110000011110011100;
            12'b010110110010: out = 32'b00000000000000110000011101001000;
            12'b010110110011: out = 32'b00000000000000110000011011110100;
            12'b010110110100: out = 32'b00000000000000110000011010100001;
            12'b010110110101: out = 32'b00000000000000110000011001001101;
            12'b010110110110: out = 32'b00000000000000110000010111111001;
            12'b010110110111: out = 32'b00000000000000110000010110100101;
            12'b010110111000: out = 32'b00000000000000110000010101010010;
            12'b010110111001: out = 32'b00000000000000110000010011111110;
            12'b010110111010: out = 32'b00000000000000110000010010101010;
            12'b010110111011: out = 32'b00000000000000110000010001010110;
            12'b010110111100: out = 32'b00000000000000110000010000000010;
            12'b010110111101: out = 32'b00000000000000110000001110101101;
            12'b010110111110: out = 32'b00000000000000110000001101011001;
            12'b010110111111: out = 32'b00000000000000110000001100000101;
            12'b010111000000: out = 32'b00000000000000110000001010110001;
            12'b010111000001: out = 32'b00000000000000110000001001011100;
            12'b010111000010: out = 32'b00000000000000110000001000001000;
            12'b010111000011: out = 32'b00000000000000110000000110110100;
            12'b010111000100: out = 32'b00000000000000110000000101011111;
            12'b010111000101: out = 32'b00000000000000110000000100001011;
            12'b010111000110: out = 32'b00000000000000110000000010110110;
            12'b010111000111: out = 32'b00000000000000110000000001100010;
            12'b010111001000: out = 32'b00000000000000110000000000001101;
            12'b010111001001: out = 32'b00000000000000101111111110111000;
            12'b010111001010: out = 32'b00000000000000101111111101100100;
            12'b010111001011: out = 32'b00000000000000101111111100001111;
            12'b010111001100: out = 32'b00000000000000101111111010111010;
            12'b010111001101: out = 32'b00000000000000101111111001100101;
            12'b010111001110: out = 32'b00000000000000101111111000010000;
            12'b010111001111: out = 32'b00000000000000101111110110111011;
            12'b010111010000: out = 32'b00000000000000101111110101100110;
            12'b010111010001: out = 32'b00000000000000101111110100010001;
            12'b010111010010: out = 32'b00000000000000101111110010111100;
            12'b010111010011: out = 32'b00000000000000101111110001100111;
            12'b010111010100: out = 32'b00000000000000101111110000010010;
            12'b010111010101: out = 32'b00000000000000101111101110111101;
            12'b010111010110: out = 32'b00000000000000101111101101100111;
            12'b010111010111: out = 32'b00000000000000101111101100010010;
            12'b010111011000: out = 32'b00000000000000101111101010111101;
            12'b010111011001: out = 32'b00000000000000101111101001100111;
            12'b010111011010: out = 32'b00000000000000101111101000010010;
            12'b010111011011: out = 32'b00000000000000101111100110111100;
            12'b010111011100: out = 32'b00000000000000101111100101100111;
            12'b010111011101: out = 32'b00000000000000101111100100010001;
            12'b010111011110: out = 32'b00000000000000101111100010111011;
            12'b010111011111: out = 32'b00000000000000101111100001100110;
            12'b010111100000: out = 32'b00000000000000101111100000010000;
            12'b010111100001: out = 32'b00000000000000101111011110111010;
            12'b010111100010: out = 32'b00000000000000101111011101100100;
            12'b010111100011: out = 32'b00000000000000101111011100001110;
            12'b010111100100: out = 32'b00000000000000101111011010111000;
            12'b010111100101: out = 32'b00000000000000101111011001100010;
            12'b010111100110: out = 32'b00000000000000101111011000001100;
            12'b010111100111: out = 32'b00000000000000101111010110110110;
            12'b010111101000: out = 32'b00000000000000101111010101100000;
            12'b010111101001: out = 32'b00000000000000101111010100001010;
            12'b010111101010: out = 32'b00000000000000101111010010110100;
            12'b010111101011: out = 32'b00000000000000101111010001011101;
            12'b010111101100: out = 32'b00000000000000101111010000000111;
            12'b010111101101: out = 32'b00000000000000101111001110110001;
            12'b010111101110: out = 32'b00000000000000101111001101011010;
            12'b010111101111: out = 32'b00000000000000101111001100000100;
            12'b010111110000: out = 32'b00000000000000101111001010101101;
            12'b010111110001: out = 32'b00000000000000101111001001010111;
            12'b010111110010: out = 32'b00000000000000101111001000000000;
            12'b010111110011: out = 32'b00000000000000101111000110101010;
            12'b010111110100: out = 32'b00000000000000101111000101010011;
            12'b010111110101: out = 32'b00000000000000101111000011111100;
            12'b010111110110: out = 32'b00000000000000101111000010100110;
            12'b010111110111: out = 32'b00000000000000101111000001001111;
            12'b010111111000: out = 32'b00000000000000101110111111111000;
            12'b010111111001: out = 32'b00000000000000101110111110100001;
            12'b010111111010: out = 32'b00000000000000101110111101001010;
            12'b010111111011: out = 32'b00000000000000101110111011110011;
            12'b010111111100: out = 32'b00000000000000101110111010011100;
            12'b010111111101: out = 32'b00000000000000101110111001000101;
            12'b010111111110: out = 32'b00000000000000101110110111101110;
            12'b010111111111: out = 32'b00000000000000101110110110010111;
            12'b011000000000: out = 32'b00000000000000101110110100111111;
            12'b011000000001: out = 32'b00000000000000101110110011101000;
            12'b011000000010: out = 32'b00000000000000101110110010010001;
            12'b011000000011: out = 32'b00000000000000101110110000111001;
            12'b011000000100: out = 32'b00000000000000101110101111100010;
            12'b011000000101: out = 32'b00000000000000101110101110001011;
            12'b011000000110: out = 32'b00000000000000101110101100110011;
            12'b011000000111: out = 32'b00000000000000101110101011011011;
            12'b011000001000: out = 32'b00000000000000101110101010000100;
            12'b011000001001: out = 32'b00000000000000101110101000101100;
            12'b011000001010: out = 32'b00000000000000101110100111010101;
            12'b011000001011: out = 32'b00000000000000101110100101111101;
            12'b011000001100: out = 32'b00000000000000101110100100100101;
            12'b011000001101: out = 32'b00000000000000101110100011001101;
            12'b011000001110: out = 32'b00000000000000101110100001110101;
            12'b011000001111: out = 32'b00000000000000101110100000011101;
            12'b011000010000: out = 32'b00000000000000101110011111000110;
            12'b011000010001: out = 32'b00000000000000101110011101101110;
            12'b011000010010: out = 32'b00000000000000101110011100010101;
            12'b011000010011: out = 32'b00000000000000101110011010111101;
            12'b011000010100: out = 32'b00000000000000101110011001100101;
            12'b011000010101: out = 32'b00000000000000101110011000001101;
            12'b011000010110: out = 32'b00000000000000101110010110110101;
            12'b011000010111: out = 32'b00000000000000101110010101011101;
            12'b011000011000: out = 32'b00000000000000101110010100000100;
            12'b011000011001: out = 32'b00000000000000101110010010101100;
            12'b011000011010: out = 32'b00000000000000101110010001010011;
            12'b011000011011: out = 32'b00000000000000101110001111111011;
            12'b011000011100: out = 32'b00000000000000101110001110100011;
            12'b011000011101: out = 32'b00000000000000101110001101001010;
            12'b011000011110: out = 32'b00000000000000101110001011110001;
            12'b011000011111: out = 32'b00000000000000101110001010011001;
            12'b011000100000: out = 32'b00000000000000101110001001000000;
            12'b011000100001: out = 32'b00000000000000101110000111100111;
            12'b011000100010: out = 32'b00000000000000101110000110001111;
            12'b011000100011: out = 32'b00000000000000101110000100110110;
            12'b011000100100: out = 32'b00000000000000101110000011011101;
            12'b011000100101: out = 32'b00000000000000101110000010000100;
            12'b011000100110: out = 32'b00000000000000101110000000101011;
            12'b011000100111: out = 32'b00000000000000101101111111010010;
            12'b011000101000: out = 32'b00000000000000101101111101111001;
            12'b011000101001: out = 32'b00000000000000101101111100100000;
            12'b011000101010: out = 32'b00000000000000101101111011000111;
            12'b011000101011: out = 32'b00000000000000101101111001101110;
            12'b011000101100: out = 32'b00000000000000101101111000010100;
            12'b011000101101: out = 32'b00000000000000101101110110111011;
            12'b011000101110: out = 32'b00000000000000101101110101100010;
            12'b011000101111: out = 32'b00000000000000101101110100001000;
            12'b011000110000: out = 32'b00000000000000101101110010101111;
            12'b011000110001: out = 32'b00000000000000101101110001010110;
            12'b011000110010: out = 32'b00000000000000101101101111111100;
            12'b011000110011: out = 32'b00000000000000101101101110100011;
            12'b011000110100: out = 32'b00000000000000101101101101001001;
            12'b011000110101: out = 32'b00000000000000101101101011101111;
            12'b011000110110: out = 32'b00000000000000101101101010010110;
            12'b011000110111: out = 32'b00000000000000101101101000111100;
            12'b011000111000: out = 32'b00000000000000101101100111100010;
            12'b011000111001: out = 32'b00000000000000101101100110001000;
            12'b011000111010: out = 32'b00000000000000101101100100101111;
            12'b011000111011: out = 32'b00000000000000101101100011010101;
            12'b011000111100: out = 32'b00000000000000101101100001111011;
            12'b011000111101: out = 32'b00000000000000101101100000100001;
            12'b011000111110: out = 32'b00000000000000101101011111000111;
            12'b011000111111: out = 32'b00000000000000101101011101101101;
            12'b011001000000: out = 32'b00000000000000101101011100010011;
            12'b011001000001: out = 32'b00000000000000101101011010111000;
            12'b011001000010: out = 32'b00000000000000101101011001011110;
            12'b011001000011: out = 32'b00000000000000101101011000000100;
            12'b011001000100: out = 32'b00000000000000101101010110101010;
            12'b011001000101: out = 32'b00000000000000101101010101001111;
            12'b011001000110: out = 32'b00000000000000101101010011110101;
            12'b011001000111: out = 32'b00000000000000101101010010011011;
            12'b011001001000: out = 32'b00000000000000101101010001000000;
            default: out = 0;
        endcase
    end

endmodule: cossine_lut
