module cossine_lut
(
    input logic [31:0]in,
    output logic [31:0]out
);

endmodule: cossine_lut
