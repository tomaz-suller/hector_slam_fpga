`ifndef HSLAM

`define HSLAM
`define VSIZE 32

`endif
