`include "../packages.sv"

module cossine_lut
    import fixed_pkg::fixed_t;
(
    input fixed_t in,
    output fixed_t out
);

endmodule: cossine_lut
